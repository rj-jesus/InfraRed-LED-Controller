library IEEE;
use IEEE.STD_LOGIC_1164.all;
--use IEEE.NUMERIC_STD.all;

entity SoundRom is
  port(iClk   : in std_logic;
       iRst   : in std_logic;
       iEn    : in std_logic;
       oDataL : out std_logic_vector(15 downto 0);
       oDataR : out std_logic_vector(15 downto 0));
end SoundRom;

architecture RTL of SoundRom is
  constant ArraySize : natural := 81648;
  type TROM is array(0 to ArraySize-1) of std_logic_vector(15 downto 0);
  constant SoundL : TROM := (x"09F7", x"0AB1", x"09A2", x"0A6E", x"0954", x"09CF", x"090C", x"091A", x"08C4", x"086B", x"085A", x"07E9", x"07FC", x"077D", x"0775", x"0710", x"06E1", x"069E", x"064E", x"062C", x"05C4", x"059F", x"0532", x"04FF", x"049E", x"0444", x"03EB", x"037F", x"0340", x"02E5", x"02C1", x"0280", x"0252", x"0210", x"01C2", x"017A", x"0122", x"00E4", x"008B", x"004B", x"0001", x"FFC8", x"FF89", x"FF43", x"FF02", x"FEB0", x"FE7D", x"FE3B", x"FE0E", x"FDD1", x"FD9E", x"FD68", x"FD34", x"FD02", x"FCD0", x"FCA4", x"FC73", x"FC47", x"FC19", x"FBEB", x"FBBA", x"FB7D", x"FB35", x"FAE9", x"FA92", x"FA49", x"F9F4", x"F9AA", x"F955", x"F90B", x"F8BA", x"F878", x"F833", x"F7F4", x"F7BB", x"F77E", x"F750", x"F720", x"F6F9", x"F6C4", x"F68E", x"F652", x"F615", x"F5E0", x"F5AE", x"F57D", x"F54D", x"F50C", x"F4CC", x"F480", x"F432", x"F3E3", x"F391", x"F343", x"F2F7", x"F2A3", x"F24F", x"F1F7", x"F1A7", x"F165", x"F11D", x"F0DD", x"F09C", x"F061", x"F02F", x"EFF6", x"EFA5", x"EF49", x"EEDC", x"EE84", x"EE36", x"EDF4", x"EDB5", x"ED6A", x"ED20", x"ECDA", x"EC97", x"EC62", x"EC25", x"EBF0", x"EBB4", x"EB89", x"EB5C", x"EB38", x"EB14", x"EADA", x"EAA0", x"EA4E", x"EA10", x"E9D4", x"E9B4", x"E98E", x"E967", x"E932", x"E8F3", x"E8B5", x"E87F", x"E84C", x"E81E", x"E7EC", x"E7BA", x"E782", x"E75B", x"E741", x"E716", x"E6F0", x"E6CB", x"E6B8", x"E696", x"E671", x"E654", x"E62B", x"E600", x"E5CF", x"E5C0", x"E5B1", x"E5B9", x"E5A3", x"E591", x"E564", x"E547", x"E525", x"E508", x"E4EC", x"E4CB", x"E4AB", x"E489", x"E471", x"E455", x"E449", x"E430", x"E417", x"E3EE", x"E3CB", x"E3BC", x"E3BE", x"E3CE", x"E3D7", x"E3D5", x"E3C2", x"E3B3", x"E3A0", x"E393", x"E380", x"E363", x"E341", x"E322", x"E303", x"E2EE", x"E2DA", x"E2C3", x"E2A1", x"E286", x"E263", x"E252", x"E23C", x"E230", x"E213", x"E201", x"E1EA", x"E1DF", x"E1CC", x"E1BF", x"E1A4", x"E193", x"E17D", x"E175", x"E16F", x"E16C", x"E16B", x"E165", x"E162", x"E156", x"E14A", x"E13A", x"E125", x"E100", x"E0DB", x"E0C3", x"E0AD", x"E0B2", x"E0BA", x"E0C5", x"E0C6", x"E0D1", x"E0DF", x"E0EE", x"E0FC", x"E106", x"E111", x"E11E", x"E132", x"E141", x"E152", x"E14E", x"E151", x"E14F", x"E156", x"E16C", x"E17D", x"E19D", x"E1AF", x"E1CC", x"E1E1", x"E1F5", x"E209", x"E209", x"E21A", x"E21F", x"E23D", x"E264", x"E29A", x"E2CD", x"E2FE", x"E317", x"E331", x"E340", x"E35A", x"E371", x"E37A", x"E373", x"E363", x"E35A", x"E36B", x"E396", x"E3C7", x"E3F6", x"E414", x"E435", x"E457", x"E491", x"E4C0", x"E4E5", x"E4F3", x"E4F9", x"E500", x"E521", x"E53D", x"E55C", x"E567", x"E56B", x"E56A", x"E56D", x"E57C", x"E597", x"E5AE", x"E5BE", x"E5D8", x"E5EC", x"E60D", x"E61B", x"E625", x"E61C", x"E617", x"E620", x"E643", x"E67F", x"E6AA", x"E6D1", x"E6D4", x"E6DD", x"E6E7", x"E6FC", x"E71A", x"E72A", x"E734", x"E731", x"E73E", x"E765", x"E7A5", x"E7F7", x"E83E", x"E874", x"E88E", x"E8A4", x"E8BC", x"E8D3", x"E8EA", x"E8FD", x"E904", x"E905", x"E911", x"E922", x"E943", x"E960", x"E97A", x"E98D", x"E994", x"E9A9", x"E9D6", x"EA06", x"EA4D", x"EA84", x"EAB6", x"EAE1", x"EAFD", x"EB20", x"EB2B", x"EB37", x"EB43", x"EB53", x"EB71", x"EB90", x"EBBA", x"EBD8", x"EC01", x"EC27", x"EC54", x"EC7D", x"ECB5", x"ECE2", x"ED0C", x"ED26", x"ED48", x"ED6E", x"ED9B", x"EDC7", x"EDD5", x"EDD2", x"EDB6", x"ED9F", x"ED91", x"ED9C", x"EDBA", x"EDDF", x"EE02", x"EE0F", x"EE16", x"EE1E", x"EE25", x"EE41", x"EE5A", x"EE67", x"EE6E", x"EE6C", x"EE6E", x"EE6C", x"EE6E", x"EE77", x"EE77", x"EE79", x"EE8E", x"EE9B", x"EEA8", x"EEBC", x"EECE", x"EECC", x"EED6", x"EEE1", x"EEF1", x"EF08", x"EF25", x"EF3E", x"EF44", x"EF61", x"EF6C", x"EF7D", x"EF7D", x"EF82", x"EF7C", x"EF80", x"EF8F", x"EF94", x"EF9F", x"EFA9", x"EFB3", x"EFBF", x"EFDE", x"EFFB", x"F025", x"F04F", x"F074", x"F06E", x"F06E", x"F073", x"F077", x"F09D", x"F0CB", x"F0F7", x"F108", x"F12B", x"F142", x"F155", x"F194", x"F1D1", x"F1E9", x"F203", x"F22A", x"F24F", x"F253", x"F272", x"F27F", x"F282", x"F294", x"F2A7", x"F2B5", x"F2C3", x"F2D3", x"F2CD", x"F2D0", x"F2DE", x"F2F5", x"F30D", x"F335", x"F354", x"F365", x"F382", x"F3A4", x"F3C0", x"F3E2", x"F404", x"F40D", x"F412", x"F439", x"F454", x"F481", x"F4AD", x"F4CD", x"F4BC", x"F4B6", x"F4BF", x"F4C0", x"F4E0", x"F511", x"F533", x"F545", x"F54F", x"F54F", x"F538", x"F52C", x"F531", x"F543", x"F55F", x"F574", x"F587", x"F589", x"F59C", x"F5B5", x"F5EC", x"F61B", x"F63D", x"F652", x"F66E", x"F66C", x"F67C", x"F699", x"F6C6", x"F6F1", x"F72F", x"F768", x"F773", x"F778", x"F792", x"F79A", x"F7B3", x"F7DB", x"F7FF", x"F804", x"F81B", x"F845", x"F86B", x"F895", x"F8C8", x"F8E1", x"F8EF", x"F913", x"F948", x"F979", x"F9AD", x"F9EA", x"FA0F", x"FA27", x"FA27", x"FA24", x"FA2C", x"FA48", x"FA9D", x"FAF9", x"FB70", x"FBC3", x"FC1A", x"FC6A", x"FCAF", x"FCF1", x"FD38", x"FD73", x"FD93", x"FDC4", x"FDFB", x"FE1D", x"FE36", x"FE68", x"FE9C", x"FEBD", x"FEEE", x"FF14", x"FF13", x"FF1C", x"FF60", x"FFB9", x"000F", x"006C", x"00B6", x"00C3", x"00D6", x"010F", x"0137", x"0158", x"018E", x"01BC", x"01E7", x"0226", x"027C", x"02B0", x"02D8", x"02FF", x"0312", x"0320", x"0355", x"038B", x"03C5", x"0413", x"0471", x"04B1", x"04F0", x"052A", x"053C", x"054E", x"055F", x"0573", x"058A", x"05BB", x"05F4", x"0614", x"064A", x"067A", x"06AA", x"06EC", x"073B", x"0774", x"079E", x"07C5", x"07F0", x"0820", x"087C", x"08D1", x"0908", x"0939", x"0957", x"0965", x"0989", x"09C9", x"0A10", x"0A60", x"0AC1", x"0B12", x"0B62", x"0BB0", x"0BF9", x"0C25", x"0C5B", x"0C8D", x"0CBA", x"0CFA", x"0D43", x"0D76", x"0DAA", x"0DDD", x"0E02", x"0E2D", x"0E6E", x"0ED2", x"0F2F", x"0FAE", x"1024", x"1094", x"1112", x"117E", x"11D9", x"121C", x"1263", x"1291", x"12D3", x"1310", x"1337", x"1352", x"1368", x"1382", x"138D", x"13C0", x"1407", x"144C", x"1497", x"14E5", x"1518", x"154D", x"1598", x"15F2", x"164D", x"16AD", x"1700", x"172A", x"1762", x"1789", x"17B3", x"17CE", x"17F6", x"1818", x"1842", x"186A", x"1889", x"188E", x"189B", x"18B0", x"18C8", x"18F4", x"1924", x"1962", x"199D", x"19DE", x"1A03", x"1A28", x"1A3C", x"1A56", x"1A5C", x"1A82", x"1AA0", x"1AD2", x"1B0A", x"1B48", x"1B7B", x"1B8A", x"1BA3", x"1BC7", x"1BEB", x"1C1C", x"1C5F", x"1C86", x"1C8C", x"1C8D", x"1C9A", x"1C96", x"1CA4", x"1CCF", x"1CF1", x"1D07", x"1D49", x"1D90", x"1DB8", x"1DE4", x"1E06", x"1E1E", x"1E4C", x"1EA0", x"1EEB", x"1F11", x"1F34", x"1F61", x"1F89", x"1FC9", x"201B", x"2049", x"2072", x"2090", x"20B2", x"20BC", x"20DA", x"20E0", x"20D4", x"20D8", x"20C5", x"20C6", x"20C7", x"20DF", x"20D0", x"20C3", x"20AB", x"2086", x"206F", x"2092", x"20B4", x"20D0", x"20EF", x"2100", x"20F3", x"2102", x"212F", x"2155", x"2174", x"21AB", x"21CC", x"21E7", x"2206", x"220D", x"21F3", x"21D2", x"21A9", x"2193", x"2174", x"2173", x"215B", x"214D", x"213F", x"211A", x"20FE", x"20E8", x"20C4", x"20A4", x"208D", x"2059", x"2018", x"1FF1", x"1FDE", x"1FCE", x"1FD2", x"1FED", x"1FE7", x"1FF3", x"2016", x"2035", x"202B", x"202C", x"2019", x"1FF2", x"1FF0", x"1FFF", x"2004", x"1FE8", x"1FC9", x"1F82", x"1F3F", x"1F10", x"1EF4", x"1ED4", x"1EB7", x"1E89", x"1E47", x"1E07", x"1DC5", x"1D85", x"1D68", x"1D58", x"1D37", x"1D24", x"1D27", x"1D1D", x"1D24", x"1D42", x"1D42", x"1D19", x"1D1A", x"1D30", x"1D3E", x"1D41", x"1D4F", x"1D24", x"1CEC", x"1CE5", x"1CEB", x"1CCF", x"1CBA", x"1CB3", x"1C89", x"1C61", x"1C4C", x"1C19", x"1BCF", x"1B99", x"1B73", x"1B4F", x"1B43", x"1B40", x"1B2D", x"1B00", x"1AD7", x"1AAA", x"1A81", x"1A68", x"1A54", x"1A2A", x"19F6", x"19B8", x"196C", x"1917", x"18D8", x"18A5", x"1885", x"1878", x"185F", x"1845", x"181A", x"17E9", x"17A8", x"1759", x"1710", x"16C8", x"168B", x"1661", x"1632", x"15EF", x"15B2", x"1580", x"1543", x"1505", x"14D2", x"14A7", x"1486", x"147E", x"147D", x"1467", x"142E", x"140E", x"13EC", x"13CB", x"13BE", x"13A6", x"136C", x"1319", x"12BD", x"1258", x"11F5", x"11A3", x"115D", x"1127", x"10FD", x"10CC", x"10A5", x"1081", x"107A", x"1083", x"10B0", x"10D0", x"10E8", x"10FB", x"1105", x"10F4", x"10D1", x"1099", x"1049", x"0FFB", x"0FD9", x"0FAE", x"0F87", x"0F6B", x"0F37", x"0F08", x"0EDF", x"0EC4", x"0E98", x"0E7B", x"0E6D", x"0E73", x"0E6F", x"0E82", x"0E7B", x"0E45", x"0E0A", x"0DC2", x"0D7F", x"0D5A", x"0D59", x"0D45", x"0D2A", x"0CFA", x"0CBD", x"0C7C", x"0C5D", x"0C51", x"0C3F", x"0C3D", x"0C1F", x"0BF1", x"0BC8", x"0BAE", x"0B8F", x"0B72", x"0B4D", x"0AF2", x"0A88", x"0A2F", x"09E4", x"09A2", x"0988", x"0970", x"0950", x"094A", x"0950", x"092F", x"0900", x"08C8", x"0885", x"0837", x"081D", x"0805", x"07D7", x"07CE", x"07BC", x"0796", x"0774", x"0772", x"0741", x"06FE", x"06C8", x"069B", x"066C", x"0683", x"06B8", x"06A0", x"0664", x"0615", x"05BE", x"0561", x"053E", x"0523", x"04ED", x"04B9", x"049A", x"0472", x"043D", x"0420", x"040A", x"03FA", x"03F7", x"03F5", x"03F2", x"03F6", x"041B", x"0450", x"0489", x"04A9", x"04AD", x"0486", x"044D", x"03FB", x"03B4", x"0377", x"0351", x"0347", x"0352", x"0355", x"0339", x"0323", x"02E8", x"02B7", x"0294", x"029E", x"027B", x"024E", x"021C", x"01EC", x"01B5", x"01B0", x"01A0", x"015B", x"0100", x"00CD", x"00A3", x"009B", x"00B0", x"00C7", x"00B7", x"0098", x"0086", x"0058", x"003D", x"002F", x"002F", x"0031", x"0036", x"0021", x"000D", x"0000", x"FFEF", x"FFC3", x"FFA6", x"FF72", x"FF1F", x"FEE4", x"FEAC", x"FE5C", x"FE12", x"FE00", x"FDF2", x"FDEF", x"FDFE", x"FDE1", x"FD81", x"FD2D", x"FD06", x"FCE6", x"FD0B", x"FD3A", x"FD36", x"FCFA", x"FCD8", x"FCA6", x"FC7D", x"FC80", x"FC7C", x"FC40", x"FC0F", x"FBF8", x"FBCD", x"FBC0", x"FBC6", x"FB9E", x"FB49", x"FB1A", x"FAD5", x"FA96", x"FA95", x"FA8C", x"FA4B", x"FA16", x"F9EF", x"F9AA", x"F983", x"F997", x"F97B", x"F93C", x"F93D", x"F947", x"F924", x"F935", x"F93F", x"F8FD", x"F8BF", x"F8CD", x"F8CD", x"F8BA", x"F8C0", x"F894", x"F81F", x"F7D1", x"F7C7", x"F7B8", x"F7BF", x"F7D1", x"F7A2", x"F75A", x"F715", x"F6D8", x"F6AB", x"F690", x"F66E", x"F627", x"F5D7", x"F57F", x"F51D", x"F4F5", x"F4D6", x"F4AB", x"F480", x"F46F", x"F438", x"F41A", x"F412", x"F3E1", x"F395", x"F354", x"F314", x"F2CE", x"F2B2", x"F2AC", x"F26A", x"F22D", x"F1F1", x"F1B0", x"F175", x"F166", x"F12F", x"F0CE", x"F085", x"F048", x"F01B", x"F003", x"EFF5", x"EFB8", x"EF67", x"EF24", x"EEEE", x"EEC2", x"EEA4", x"EE64", x"EE15", x"EDA8", x"ED38", x"ECD4", x"ECB2", x"EC98", x"EC88", x"EC7F", x"EC67", x"EC2B", x"EC15", x"EC1F", x"EC23", x"EC2D", x"EC3B", x"EC1E", x"EBE7", x"EBD4", x"EBB3", x"EB9F", x"EB8E", x"EB7A", x"EB2A", x"EAEA", x"EAB9", x"EA73", x"EA37", x"EA1E", x"E9F6", x"E9E4", x"E9FB", x"EA1E", x"E9FC", x"E9D9", x"E99D", x"E958", x"E91B", x"E8FD", x"E8CB", x"E89D", x"E872", x"E83D", x"E810", x"E7DE", x"E79A", x"E75D", x"E735", x"E700", x"E6C8", x"E6C1", x"E6CC", x"E6E4", x"E714", x"E736", x"E6FB", x"E6A7", x"E66E", x"E626", x"E603", x"E608", x"E5F0", x"E5A0", x"E57C", x"E56F", x"E561", x"E582", x"E5A9", x"E564", x"E4FA", x"E488", x"E40A", x"E3A0", x"E386", x"E37C", x"E33F", x"E327", x"E315", x"E2DE", x"E2BA", x"E2A8", x"E25B", x"E1FD", x"E1C5", x"E182", x"E144", x"E13A", x"E121", x"E0CF", x"E08D", x"E05E", x"E024", x"E012", x"E03C", x"E039", x"E02A", x"E059", x"E084", x"E093", x"E0A8", x"E087", x"E01C", x"DFBC", x"DFA7", x"DF96", x"DF90", x"DFA5", x"DF8F", x"DF65", x"DF69", x"DFA0", x"DFCA", x"E013", x"E037", x"E028", x"DFFB", x"DFDD", x"DFCD", x"DFD6", x"DFFB", x"E017", x"E014", x"E026", x"E041", x"E047", x"E05D", x"E064", x"E040", x"E00D", x"DFFA", x"DFF3", x"DFE6", x"E000", x"E019", x"E032", x"E050", x"E093", x"E0C8", x"E0E3", x"E10C", x"E13D", x"E162", x"E18F", x"E1A8", x"E18C", x"E146", x"E104", x"E0DE", x"E0BA", x"E0C5", x"E0D5", x"E0DB", x"E0DF", x"E108", x"E12E", x"E155", x"E187", x"E1B1", x"E1B6", x"E1B1", x"E1BC", x"E1AB", x"E19E", x"E19C", x"E189", x"E175", x"E170", x"E178", x"E188", x"E1A5", x"E1B7", x"E1B7", x"E1B7", x"E1C7", x"E1B7", x"E1CF", x"E1E9", x"E1EE", x"E1F6", x"E21D", x"E244", x"E254", x"E271", x"E29E", x"E2AC", x"E2FA", x"E373", x"E3E1", x"E41B", x"E44B", x"E446", x"E42E", x"E43C", x"E45D", x"E46D", x"E495", x"E4C7", x"E4EF", x"E521", x"E570", x"E59B", x"E5B6", x"E5E2", x"E5F9", x"E608", x"E64C", x"E6A0", x"E6E3", x"E72E", x"E760", x"E75F", x"E755", x"E77D", x"E7A8", x"E7EA", x"E856", x"E8AA", x"E8E5", x"E938", x"E9A0", x"E9CC", x"EA09", x"EA3D", x"EA3C", x"EA3C", x"EA64", x"EA7E", x"EA73", x"EA86", x"EAAB", x"EAC0", x"EB1B", x"EB8C", x"EBDF", x"EC16", x"EC61", x"EC8A", x"ECBE", x"ED2F", x"EDA8", x"EE10", x"EE84", x"EEF2", x"EF1F", x"EF58", x"EFA6", x"EFBC", x"EFBE", x"EFD4", x"EFD8", x"EFD3", x"F004", x"F04C", x"F050", x"F052", x"F05D", x"F058", x"F06F", x"F0D0", x"F141", x"F18D", x"F1F0", x"F249", x"F280", x"F2AF", x"F2DF", x"F2DB", x"F2C3", x"F2C3", x"F2E5", x"F30A", x"F344", x"F379", x"F38F", x"F3BF", x"F3FE", x"F457", x"F4B9", x"F518", x"F568", x"F5A7", x"F5DC", x"F5F9", x"F613", x"F644", x"F680", x"F6B3", x"F6F5", x"F72B", x"F744", x"F767", x"F79F", x"F7B8", x"F7C7", x"F7F5", x"F819", x"F842", x"F875", x"F8A6", x"F8A1", x"F8AB", x"F8D6", x"F924", x"F975", x"F9DF", x"FA36", x"FA74", x"FABB", x"FB2C", x"FB95", x"FBF5", x"FC52", x"FCB3", x"FD15", x"FD70", x"FDDB", x"FE26", x"FE52", x"FE78", x"FEA8", x"FED1", x"FEDE", x"FEF9", x"FF15", x"FF29", x"FF42", x"FF5E", x"FF5E", x"FF48", x"FF61", x"FFAD", x"0002", x"0089", x"0104", x"0149", x"016E", x"0191", x"019C", x"01A9", x"01D0", x"01F9", x"0218", x"024A", x"0284", x"029A", x"02A8", x"02C3", x"02C9", x"02E5", x"0316", x"033A", x"0347", x"0361", x"0367", x"0361", x"038B", x"03BA", x"03EA", x"041E", x"0451", x"0437", x"041D", x"042A", x"0435", x"0440", x"046D", x"0487", x"0473", x"0487", x"04C0", x"04D2", x"04E0", x"04F6", x"04E1", x"04CD", x"04F4", x"0537", x"057E", x"05EC", x"0641", x"0668", x"0694", x"06D2", x"0705", x"075C", x"07CB", x"081D", x"084D", x"08A4", x"08D2", x"08E4", x"08F9", x"0900", x"08D2", x"08D7", x"0903", x"090E", x"0925", x"0935", x"090F", x"08EA", x"091F", x"096D", x"09B4", x"0A21", x"0A6C", x"0A63", x"0A7C", x"0ACB", x"0AEC", x"0B2A", x"0B87", x"0BCB", x"0BE7", x"0C49", x"0C9F", x"0CBF", x"0CE1", x"0CE5", x"0C96", x"0C55", x"0C4A", x"0C43", x"0C4D", x"0C92", x"0CB3", x"0CBA", x"0CFB", x"0D44", x"0D65", x"0D9F", x"0DD2", x"0DCD", x"0DCE", x"0E02", x"0E15", x"0E07", x"0E15", x"0DED", x"0DB6", x"0DB2", x"0DDA", x"0DEA", x"0E0F", x"0E28", x"0E16", x"0E14", x"0E47", x"0E70", x"0E85", x"0EAB", x"0E96", x"0E49", x"0E1B", x"0E0E", x"0DE4", x"0DF7", x"0E22", x"0E2F", x"0E3B", x"0E8B", x"0EC9", x"0ED1", x"0EE2", x"0EC5", x"0E84", x"0E66", x"0E90", x"0E9E", x"0EA3", x"0EBA", x"0ECC", x"0EC5", x"0EDA", x"0EEA", x"0EBB", x"0E86", x"0E83", x"0E8D", x"0EB8", x"0F04", x"0F46", x"0F5F", x"0F7F", x"0FA2", x"0FD6", x"100D", x"1061", x"10AF", x"10F9", x"112E", x"114A", x"113E", x"111E", x"10EF", x"10E5", x"10D8", x"10CB", x"10B8", x"10AD", x"10AE", x"10B6", x"10E9", x"1128", x"115A", x"11B7", x"1240", x"12C3", x"1324", x"1382", x"13C8", x"13E8", x"141D", x"1466", x"1491", x"1494", x"14CE", x"1509", x"154E", x"159E", x"15F1", x"1612", x"1615", x"163A", x"165F", x"167E", x"16A7", x"16B1", x"1698", x"1675", x"165F", x"1653", x"1654", x"167A", x"1692", x"16C1", x"16DC", x"16F2", x"16EB", x"16E6", x"16E8", x"16F6", x"1703", x"16F3", x"16D5", x"16BE", x"16A5", x"1683", x"1686", x"168C", x"1688", x"16CB", x"1748", x"1795", x"17BC", x"17EB", x"17E8", x"17C7", x"17DF", x"17F8", x"17B5", x"1772", x"1768", x"175C", x"177B", x"17F2", x"1832", x"182F", x"183B", x"1857", x"185D", x"1890", x"18CD", x"18A4", x"1845", x"17F7", x"1796", x"1744", x"1755", x"178A", x"17AB", x"1802", x"1862", x"18AE", x"1903", x"1971", x"19A9", x"19D5", x"1A08", x"1A17", x"1A2B", x"1A71", x"1A98", x"1A95", x"1AA3", x"1AA0", x"1A6F", x"1A94", x"1AE8", x"1B09", x"1B35", x"1B89", x"1BBA", x"1BCF", x"1C15", x"1C1F", x"1BBA", x"1B80", x"1B66", x"1B51", x"1B70", x"1BB9", x"1BB7", x"1B7E", x"1B70", x"1B45", x"1B1A", x"1B2C", x"1B40", x"1B23", x"1B19", x"1B25", x"1B1F", x"1B69", x"1BF3", x"1C5A", x"1C93", x"1CBD", x"1CA6", x"1C7A", x"1C81", x"1C79", x"1C26", x"1BD7", x"1B87", x"1B1D", x"1AF6", x"1B15", x"1B02", x"1ADE", x"1ACC", x"1AA2", x"1A86", x"1ACA", x"1B27", x"1B63", x"1B9D", x"1BBC", x"1B7B", x"1B19", x"1AB2", x"1A06", x"1959", x"1900", x"18E7", x"18F7", x"1950", x"19AB", x"19D0", x"19EB", x"1A18", x"1A2B", x"1A52", x"1A85", x"1A93", x"1A81", x"1A6A", x"1A3C", x"1A03", x"19EE", x"19D8", x"198F", x"1951", x"192D", x"1913", x"194C", x"19C1", x"1A23", x"1A4B", x"1A65", x"1A72", x"1A63", x"1A6F", x"1A76", x"1A51", x"1A0B", x"19CE", x"1994", x"1962", x"1960", x"197F", x"19AF", x"19D8", x"19FE", x"19E7", x"19A1", x"193E", x"18EF", x"189E", x"1876", x"185C", x"183C", x"17E2", x"179B", x"176C", x"1734", x"170D", x"16F1", x"16B7", x"166A", x"1651", x"1666", x"165F", x"1653", x"1649", x"1617", x"15E4", x"15CF", x"15C4", x"158E", x"156D", x"1542", x"14F8", x"149F", x"1437", x"13AD", x"132F", x"12D3", x"1289", x"125E", x"1254", x"124D", x"1239", x"1239", x"123C", x"1232", x"1252", x"1274", x"126A", x"124F", x"1210", x"1191", x"10FC", x"1096", x"1031", x"0FDF", x"0FAD", x"0F91", x"0F64", x"0F72", x"0FAB", x"0FC1", x"0F9E", x"0F58", x"0EF1", x"0E6B", x"0E2D", x"0DF4", x"0DA3", x"0D3B", x"0CEA", x"0C94", x"0C4C", x"0C1C", x"0BFA", x"0BC8", x"0BB2", x"0B9D", x"0B84", x"0B4D", x"0B0D", x"0ACE", x"0A99", x"0A5E", x"0A3D", x"0A1B", x"09E3", x"09B0", x"0991", x"096A", x"0928", x"08ED", x"08B2", x"0861", x"0826", x"080C", x"07D0", x"0774", x"0721", x"06DF", x"0697", x"0675", x"0662", x"0642", x"0619", x"0611", x"05FB", x"05CD", x"059B", x"0560", x"0527", x"0500", x"04E4", x"04C4", x"0498", x"046A", x"041B", x"03BE", x"0353", x"02E4", x"0286", x"0242", x"01F2", x"019E", x"0136", x"00BB", x"0040", x"FFD1", x"FF81", x"FF43", x"FF29", x"FF2D", x"FF2A", x"FF20", x"FF06", x"FEC7", x"FE59", x"FDE1", x"FD67", x"FCEF", x"FC8A", x"FC39", x"FBFA", x"FBB1", x"FB7E", x"FB55", x"FB2A", x"FAF7", x"FACB", x"FAB9", x"FA92", x"FA79", x"FA63", x"FA56", x"FA38", x"FA41", x"FA3D", x"FA26", x"F9EC", x"F9B9", x"F97C", x"F936", x"F901", x"F8C2", x"F87F", x"F83A", x"F808", x"F7DF", x"F7AA", x"F782", x"F740", x"F6EE", x"F69C", x"F659", x"F636", x"F639", x"F655", x"F670", x"F68A", x"F690", x"F682", x"F66A", x"F649", x"F621", x"F5E4", x"F5AF", x"F56E", x"F51F", x"F4DA", x"F48D", x"F447", x"F3EA", x"F3B1", x"F383", x"F34E", x"F31B", x"F301", x"F2F8", x"F2EA", x"F310", x"F339", x"F331", x"F307", x"F2EF", x"F2C2", x"F266", x"F229", x"F1E8", x"F177", x"F10F", x"F0EF", x"F0B2", x"F068", x"F060", x"F06B", x"F04E", x"F061", x"F089", x"F06A", x"F021", x"F006", x"EFD6", x"EF94", x"EF82", x"EF80", x"EF38", x"EEFE", x"EEE9", x"EEC6", x"EEA1", x"EE91", x"EE67", x"EE10", x"EDD2", x"ED9A", x"ED71", x"ED5C", x"ED54", x"ED15", x"ECE5", x"ECAE", x"EC80", x"EC86", x"ECC7", x"ECEC", x"ECF9", x"ED24", x"ED42", x"ED41", x"ED6C", x"ED8A", x"ED59", x"ED2D", x"ED24", x"ECFD", x"ECDE", x"ECDE", x"ECBC", x"EC6B", x"EC49", x"EC44", x"EC52", x"EC8F", x"ECDA", x"ECD2", x"ECA4", x"EC7A", x"EC52", x"EC3C", x"EC71", x"EC8F", x"EC8C", x"ECB2", x"ECEA", x"ED12", x"ED51", x"ED9B", x"ED97", x"ED87", x"EDAD", x"EDBC", x"EDA3", x"EDA1", x"ED73", x"ECF0", x"ECA5", x"ECA6", x"EC87", x"EC5E", x"EC4C", x"EC22", x"EBCC", x"EBD2", x"EBF7", x"EBE2", x"EBB6", x"EBA2", x"EB84", x"EB64", x"EB73", x"EB91", x"EB87", x"EB83", x"EB87", x"EB83", x"EB7A", x"EB87", x"EBA3", x"EBD5", x"EBC6", x"EB75", x"EAEF", x"EA4D", x"E9B7", x"E999", x"E9CB", x"E9FD", x"EA04", x"EA16", x"EA00", x"E9D7", x"EA03", x"EA58", x"EA79", x"EA98", x"EACA", x"EAC2", x"EA83", x"EA4B", x"EA09", x"E989", x"E942", x"E90D", x"E8C9", x"E881", x"E88A", x"E8B9", x"E91C", x"E9A7", x"EA08", x"EA17", x"E9F5", x"E9A7", x"E944", x"E908", x"E8FC", x"E8F7", x"E91E", x"E961", x"E97C", x"E979", x"E9AC", x"E9D1", x"E9E2", x"EA04", x"EA00", x"E9B4", x"E96A", x"E979", x"E9A7", x"E9E2", x"EA30", x"EA30", x"E9CD", x"E952", x"E907", x"E8E3", x"E8EB", x"E923", x"E948", x"E934", x"E8FA", x"E8CA", x"E8DE", x"E930", x"E9CA", x"EAA1", x"EB69", x"EBE7", x"EC59", x"ECEF", x"ED6A", x"EDB7", x"EE1F", x"EE51", x"EE09", x"ED8D", x"ED08", x"EC37", x"EB76", x"EB3B", x"EB3F", x"EB0D", x"EABA", x"EA40", x"E96A", x"E8A6", x"E83B", x"E7E0", x"E76F", x"E6F0", x"E666", x"E5B8", x"E525", x"E4B0", x"E438", x"E3BB", x"E325", x"E286", x"E21B", x"E1F7", x"E238", x"E2D5", x"E384", x"E3B9", x"E374", x"E30C", x"E29A", x"E2B7", x"E3D9", x"E585", x"E705", x"E84A", x"E93A", x"E98C", x"E98A", x"E9B7", x"E99F", x"E940", x"E8FB", x"E8DE", x"E872", x"E7F5", x"E7A2", x"E73F", x"E6F9", x"E702", x"E731", x"E734", x"E728", x"E726", x"E717", x"E737", x"E782", x"E7DB", x"E82D", x"E865", x"E85D", x"E843", x"E818", x"E7CF", x"E799", x"E780", x"E757", x"E728", x"E752", x"E791", x"E79C", x"E78A", x"E72F", x"E5FB", x"E4DE", x"E4A0", x"E52D", x"E646", x"E814", x"E9C9", x"EA8E", x"EAD4", x"EADE", x"EA37", x"E921", x"E887", x"E82B", x"E7A5", x"E74A", x"E6FA", x"E64B", x"E595", x"E53C", x"E4EB", x"E485", x"E468", x"E47D", x"E4A6", x"E506", x"E577", x"E5DA", x"E656", x"E6D0", x"E724", x"E769", x"E798", x"E776", x"E75C", x"E76C", x"E748", x"E726", x"E748", x"E754", x"E70E", x"E72E", x"E749", x"E697", x"E59A", x"E4FE", x"E4A1", x"E4F7", x"E6BA", x"E8E4", x"EA54", x"EB73", x"EC96", x"ECF1", x"ECB0", x"EC95", x"EC43", x"EBBA", x"EBBD", x"EC3B", x"EC45", x"EBF6", x"EBBB", x"EB83", x"EB44", x"EB48", x"EB60", x"EB68", x"EB7E", x"EBC9", x"EC1B", x"EC6B", x"EC50", x"EBE0", x"EB46", x"EA8F", x"E9BF", x"E946", x"E91B", x"E8BE", x"E87B", x"E8A8", x"E8E5", x"E8FE", x"E9C4", x"EAE2", x"EB7C", x"EBE1", x"EC34", x"EBD2", x"EB53", x"EC64", x"EEAC", x"F119", x"F38A", x"F5B5", x"F67E", x"F666", x"F683", x"F65B", x"F57D", x"F4D1", x"F4AA", x"F461", x"F41E", x"F422", x"F3CD", x"F31C", x"F29A", x"F25B", x"F211", x"F1F1", x"F1ED", x"F1F7", x"F205", x"F230", x"F240", x"F271", x"F292", x"F26C", x"F238", x"F221", x"F1F9", x"F1E7", x"F26E", x"F2E9", x"F320", x"F39C", x"F468", x"F500", x"F5CE", x"F6C1", x"F6AE", x"F594", x"F4AB", x"F467", x"F500", x"F70C", x"FA01", x"FC43", x"FD7D", x"FE39", x"FE39", x"FD7F", x"FCD2", x"FC4F", x"FB7A", x"FAC5", x"FA53", x"F9C5", x"F93B", x"F8FF", x"F8F6", x"F8FD", x"F925", x"F957", x"F979", x"F9C6", x"F9F5", x"F9DC", x"F9C0", x"F9C2", x"F9B4", x"F9F5", x"FA7C", x"FAB2", x"FA86", x"FA8F", x"FA9F", x"FA71", x"FA95", x"FAFC", x"FB05", x"FB42", x"FC55", x"FD7F", x"FDD3", x"FDA7", x"FCFC", x"FBD8", x"FBD1", x"FDCC", x"00BE", x"0390", x"0638", x"082E", x"08F3", x"091D", x"092E", x"08B2", x"07F2", x"07A7", x"0781", x"0739", x"06DD", x"06A7", x"068F", x"06CD", x"0745", x"07CA", x"0863", x"090E", x"09B1", x"0A69", x"0AEB", x"0AC7", x"0A92", x"0ACC", x"0AF6", x"0B18", x"0B87", x"0B94", x"0AEE", x"0A94", x"0A75", x"097E", x"0870", x"081C", x"07BB", x"0726", x"073B", x"06B9", x"049B", x"029F", x"0234", x"02B4", x"0491", x"0864", x"0C06", x"0E44", x"1015", x"1180", x"118D", x"1153", x"11BB", x"11D2", x"119A", x"11FF", x"1269", x"1220", x"11F5", x"1209", x"11E3", x"11B8", x"11D7", x"119F", x"112F", x"10ED", x"10CA", x"10BD", x"10C2", x"1082", x"1010", x"100E", x"1038", x"1071", x"1138", x"120D", x"1241", x"1291", x"132F", x"132D", x"1322", x"1429", x"14FF", x"148C", x"1396", x"1200", x"0F76", x"0E0E", x"0F47", x"1189", x"13C7", x"1672", x"185B", x"1897", x"189C", x"18C7", x"17F6", x"16AA", x"15FE", x"1524", x"13E0", x"134F", x"1304", x"120A", x"1157", x"1122", x"1095", x"1015", x"102B", x"1014", x"0FA3", x"0FCF", x"104E", x"10B5", x"1174", x"1242", x"1288", x"12D1", x"13A5", x"1459", x"1507", x"15DB", x"15FE", x"158E", x"15AA", x"1631", x"16AC", x"1773", x"17EC", x"16D7", x"14E9", x"1398", x"12FD", x"1387", x"15C0", x"185D", x"19EE", x"1AD4", x"1B51", x"1B0D", x"1AC6", x"1AEF", x"1AED", x"1AA2", x"1A75", x"1A0E", x"1953", x"1903", x"18F8", x"18EF", x"193E", x"19C0", x"19CC", x"19BA", x"19AA", x"1911", x"1815", x"1747", x"168B", x"15B5", x"1561", x"1558", x"153A", x"1577", x"163E", x"1709", x"17FB", x"18F8", x"1975", x"19A2", x"1A07", x"1A96", x"1B19", x"1BA3", x"1B56", x"19D7", x"1815", x"16F8", x"16B9", x"17C2", x"19BB", x"1B61", x"1C44", x"1CD7", x"1D14", x"1D0A", x"1D6A", x"1DD4", x"1DEC", x"1DBB", x"1D5A", x"1C75", x"1B8A", x"1B06", x"1A92", x"1A50", x"1A5F", x"1A5E", x"1A37", x"1A5D", x"1A8B", x"1A7F", x"1A8D", x"1A8F", x"1A3A", x"1A14", x"1A5D", x"1A64", x"1A52", x"1A29", x"1950", x"17F7", x"1711", x"160E", x"146D", x"1317", x"1235", x"1143", x"10E7", x"111E", x"1059", x"0E5E", x"0CF7", x"0C9C", x"0D59", x"0FF4", x"13AA", x"1661", x"17D6", x"18B7", x"18AB", x"1811", x"17E9", x"17DE", x"176A", x"170A", x"16CD", x"1657", x"1613", x"161C", x"15DE", x"1574", x"1530", x"14A3", x"13E9", x"13A1", x"138C", x"13A1", x"1423", x"149E", x"14A8", x"14CD", x"151F", x"154B", x"15A1", x"15E9", x"1573", x"14EF", x"1513", x"14EC", x"146E", x"148A", x"14BA", x"14C7", x"15AC", x"16E8", x"1680", x"152F", x"1460", x"1443", x"156F", x"18FD", x"1D39", x"2057", x"2266", x"237D", x"2337", x"2285", x"221B", x"216C", x"20B9", x"203B", x"1F5B", x"1DE4", x"1C5B", x"1A78", x"187B", x"1725", x"1653", x"1597", x"159D", x"1640", x"1705", x"1835", x"19B8", x"1AB0", x"1B6D", x"1C73", x"1D0D", x"1D6B", x"1E0D", x"1DD6", x"1C74", x"1B17", x"197F", x"170F", x"14FB", x"13A1", x"1202", x"111F", x"11EA", x"129D", x"1230", x"1178", x"1054", x"0EE8", x"0F5E", x"11E4", x"14B9", x"172B", x"1915", x"1945", x"1824", x"16E6", x"1593", x"141D", x"1350", x"128E", x"1155", x"1019", x"0F21", x"0E1F", x"0DC2", x"0DF5", x"0DDF", x"0DB5", x"0DCD", x"0DAE", x"0DA0", x"0E50", x"0EFD", x"0F94", x"108C", x"1184", x"1216", x"1331", x"1490", x"1558", x"15FD", x"16C1", x"16D8", x"16C7", x"1746", x"177B", x"1774", x"183E", x"195C", x"19FB", x"1A31", x"197A", x"174B", x"151D", x"1468", x"14FB", x"16EB", x"199F", x"1B43", x"1B1D", x"19E5", x"17D6", x"1566", x"1408", x"136B", x"12C3", x"1254", x"1240", x"11D7", x"11C0", x"128B", x"1333", x"138A", x"13F2", x"13DA", x"1322", x"12AE", x"126F", x"11C4", x"1153", x"10C8", x"0F98", x"0E61", x"0DAC", x"0CBC", x"0BD9", x"0B63", x"0A81", x"093E", x"08A8", x"0833", x"0773", x"077B", x"0839", x"08DC", x"0A28", x"0BFC", x"0C74", x"0BAE", x"0B03", x"0A51", x"0A43", x"0C70", x"0FCE", x"123E", x"13ED", x"14F4", x"144C", x"1335", x"12D1", x"125D", x"1169", x"110E", x"10C6", x"1028", x"1026", x"108A", x"106E", x"100B", x"0F70", x"0DC5", x"0B9F", x"09BF", x"0794", x"0568", x"040A", x"030B", x"0246", x"029A", x"0394", x"046A", x"0580", x"06C4", x"074F", x"07BA", x"0846", x"0839", x"0806", x"088A", x"08FD", x"0991", x"0B35", x"0CAD", x"0C7F", x"0B39", x"08EF", x"0527", x"0259", x"0216", x"02C5", x"033D", x"03B4", x"02D5", x"005A", x"FE55", x"FD37", x"FBF2", x"FB0C", x"FB04", x"FAD9", x"FB26", x"FCB7", x"FEA2", x"006A", x"02B3", x"048D", x"0576", x"0667", x"0754", x"073A", x"06E4", x"06D2", x"064D", x"05E6", x"0667", x"06CE", x"0698", x"0666", x"05EE", x"04F2", x"042F", x"0382", x"023A", x"00F3", x"FFB8", x"FE24", x"FD4F", x"FDE1", x"FEB2", x"FF5C", x"FFBA", x"FE8F", x"FC29", x"FAE9", x"FB30", x"FBC3", x"FCB5", x"FD3E", x"FBB8", x"F920", x"F73B", x"F575", x"F3B0", x"F2F5", x"F2A6", x"F1B0", x"F139", x"F192", x"F19F", x"F20D", x"F396", x"F530", x"F676", x"F854", x"FA07", x"FAD0", x"FB42", x"FBCE", x"FBD2", x"FBE9", x"FC8C", x"FCE6", x"FCBA", x"FC55", x"FBBA", x"FACC", x"F9F4", x"F8F3", x"F78D", x"F622", x"F4C3", x"F38C", x"F32F", x"F37F", x"F3DF", x"F440", x"F463", x"F3B8", x"F2EC", x"F310", x"F3C8", x"F4D5", x"F656", x"F74F", x"F6DD", x"F61F", x"F57D", x"F496", x"F402", x"F454", x"F44C", x"F3FD", x"F48E", x"F594", x"F665", x"F7C9", x"F9AB", x"FAD4", x"FBA9", x"FCC1", x"FCC2", x"FB82", x"FA15", x"F897", x"F6DF", x"F5D3", x"F53B", x"F421", x"F2B1", x"F139", x"EF30", x"ED0F", x"EB4C", x"E986", x"E7F0", x"E71F", x"E6B6", x"E6AE", x"E7EE", x"E9C6", x"EAE9", x"EB6B", x"EB42", x"EA09", x"E93A", x"EA14", x"EBB8", x"EDAA", x"EFDC", x"F130", x"F123", x"F0B8", x"F010", x"EEAC", x"ED6C", x"EC43", x"EA4A", x"E84E", x"E77D", x"E6DA", x"E673", x"E6EA", x"E73A", x"E6D5", x"E721", x"E823", x"E85A", x"E828", x"E839", x"E7BE", x"E767", x"E842", x"E98D", x"EAB0", x"EC05", x"ED06", x"ED33", x"ED31", x"ECED", x"EBFA", x"EB3A", x"EAA3", x"E940", x"E7FA", x"E796", x"E6B1", x"E503", x"E364", x"E0E5", x"DD7F", x"DBB1", x"DBF4", x"DCD5", x"DE6B", x"E088", x"E177", x"E17C", x"E223", x"E2BD", x"E30C", x"E3D7", x"E471", x"E3DA", x"E360", x"E331", x"E27A", x"E20A", x"E250", x"E1FF", x"E189", x"E257", x"E36D", x"E411", x"E4E0", x"E53D", x"E42B", x"E2E0", x"E203", x"E12E", x"E106", x"E229", x"E384", x"E505", x"E6A6", x"E74C", x"E71C", x"E728", x"E67D", x"E4FC", x"E45B", x"E457", x"E3A9", x"E356", x"E30E", x"E0CA", x"DDC1", x"DCE2", x"DDA3", x"DF72", x"E340", x"E768", x"E990", x"EB2F", x"ED1B", x"EE0E", x"EE61", x"EF02", x"EECC", x"ED8C", x"ECC7", x"EC15", x"EAEB", x"EA50", x"E9FE", x"E943", x"E90E", x"E9DF", x"EA8C", x"EB3C", x"EBE5", x"EB86", x"EA6A", x"E9BC", x"E92F", x"E8DD", x"E980", x"EA73", x"EB56", x"ECA9", x"ED96", x"ED5D", x"ED39", x"ED2A", x"EC0E", x"EB2F", x"EB40", x"EAC0", x"EA2B", x"EA94", x"E958", x"E532", x"E0F0", x"DDDB", x"DBCF", x"DCFB", x"E151", x"E4E5", x"E6B4", x"E84E", x"E8AF", x"E796", x"E708", x"E6AB", x"E54A", x"E451", x"E463", x"E436", x"E441", x"E4F6", x"E506", x"E49F", x"E4E9", x"E518", x"E4F6", x"E568", x"E567", x"E3E2", x"E1FC", x"E005", x"DD87", x"DBD2", x"DBAA", x"DC13", x"DD41", x"DF87", x"E17A", x"E2EF", x"E4B1", x"E5CD", x"E606", x"E69C", x"E719", x"E70B", x"E825", x"E9F2", x"E9AD", x"E78C", x"E4DB", x"E161", x"DEF3", x"E07F", x"E456", x"E7B3", x"EAB8", x"ED59", x"EE3A", x"EEAC", x"F010", x"F10D", x"F13C", x"F1B1", x"F21B", x"F1E9", x"F1EA", x"F26E", x"F324", x"F486", x"F665", x"F7E5", x"F8EC", x"F967", x"F8E1", x"F7CC", x"F661", x"F45B", x"F201", x"EFEE", x"EE25", x"ED29", x"ED6B", x"EE52", x"EF87", x"F0DB", x"F15F", x"F0FE", x"F0C6", x"F068", x"EF4A", x"EEC6", x"EF2B", x"EEDB", x"EE33", x"ED68", x"EAB2", x"E662", x"E3DB", x"E3CB", x"E559", x"E911", x"EDB1", x"F07B", x"F19D", x"F2D0", x"F370", x"F37B", x"F458", x"F52A", x"F549", x"F5AF", x"F664", x"F671", x"F6C6", x"F78A", x"F77E", x"F703", x"F700", x"F6A1", x"F5F0", x"F618", x"F626", x"F53B", x"F461", x"F3C2", x"F2B4", x"F1F2", x"F239", x"F2D9", x"F419", x"F635", x"F818", x"F94C", x"FA06", x"F9A5", x"F850", x"F760", x"F6A7", x"F5BB", x"F56F", x"F51E", x"F324", x"F0AC", x"EF91", x"EF98", x"F141", x"F553", x"F9C6", x"FC86", x"FE4D", x"FF83", x"FF26", x"FE13", x"FD0B", x"FB79", x"F981", x"F860", x"F7EF", x"F76F", x"F738", x"F731", x"F6C6", x"F663", x"F64F", x"F64A", x"F619", x"F613", x"F641", x"F644", x"F5E6", x"F4FD", x"F384", x"F154", x"EF5C", x"EED1", x"EF47", x"EFB8", x"F074", x"F13C", x"F0EF", x"F061", x"F0D9", x"F11D", x"F09C", x"F156", x"F2C0", x"F2D9", x"F217", x"F133", x"EECD", x"EC8E", x"EDC4", x"F184", x"F5CE", x"FA99", x"FE5A", x"FEE9", x"FE1D", x"FDF1", x"FD4B", x"FC57", x"FC41", x"FBBF", x"FA81", x"FA98", x"FBFA", x"FCD3", x"FDEA", x"FF1A", x"FF1C", x"FEBE", x"FF6D", x"0034", x"00DD", x"025A", x"03C9", x"0428", x"0455", x"0410", x"02C3", x"01D3", x"016F", x"00A4", x"002C", x"0090", x"0065", x"FFB6", x"FF5E", x"FE30", x"FC34", x"FBB4", x"FC44", x"FBD9", x"FACC", x"F920", x"F5B8", x"F2A0", x"F28A", x"F47F", x"F75F", x"FB51", x"FEB8", x"FFD0", x"FFFE", x"FFF8", x"FEFF", x"FDEA", x"FD97", x"FD28", x"FCA4", x"FD36", x"FE4E", x"FF49", x"009C", x"0202", x"02A8", x"0312", x"037C", x"039B", x"03E9", x"04AD", x"0594", x"062A", x"0606", x"04BE", x"032C", x"01F2", x"00D4", x"0021", x"FFFF", x"FF62", x"FE7D", x"FE73", x"FE56", x"FD57", x"FCC3", x"FC9C", x"FBBA", x"FAD7", x"FA27", x"F7CB", x"F47C", x"F297", x"F219", x"F338", x"F742", x"FC94", x"00A8", x"0424", x"06EF", x"07C9", x"083F", x"098A", x"096D", x"07F0", x"0733", x"067B", x"058A", x"06D3", x"0901", x"0907", x"085F", x"0871", x"07C3", x"07AE", x"0A41", x"0CB8", x"0D95", x"0F28", x"10C8", x"10B0", x"10CE", x"1171", x"100D", x"0E1E", x"0DFE", x"0E14", x"0DBF", x"0E79", x"0E30", x"0BB3", x"09FA", x"09F5", x"09A7", x"096A", x"0909", x"0611", x"017A", x"FEE4", x"FE57", x"FF62", x"02EF", x"0763", x"0A53", x"0C7B", x"0E6E", x"0F0F", x"0F0B", x"0F3B", x"0EB4", x"0D97", x"0D2F", x"0D14", x"0D45", x"0EAD", x"107E", x"11B3", x"1349", x"154C", x"16DE", x"18CB", x"1B6B", x"1D17", x"1E00", x"1F45", x"2056", x"2079", x"208F", x"202D", x"1E67", x"1C5B", x"1B12", x"19FC", x"1913", x"189D", x"17F5", x"16FB", x"1660", x"1613", x"159B", x"14B2", x"12FF", x"1088", x"0E18", x"0C60", x"0BF4", x"0D72", x"1071", x"1460", x"18A4", x"1C28", x"1E17", x"1EE1", x"1F11", x"1E86", x"1E28", x"1E00", x"1CFA", x"1B63", x"1AA4", x"1A51", x"19F5", x"1A70", x"1AEC", x"19EC", x"1903", x"195E", x"198C", x"195C", x"19D7", x"19AF", x"1836", x"179F", x"1824", x"17C8", x"173F", x"1754", x"16A6", x"159E", x"1621", x"1734", x"176F", x"183E", x"19BD", x"1A6B", x"1AD5", x"1B54", x"19C6", x"1632", x"1324", x"1146", x"1097", x"123C", x"157D", x"17AE", x"18E1", x"1A38", x"1B08", x"1B13", x"1B87", x"1BC5", x"1AE9", x"1A09", x"1A00", x"1A02", x"1A12", x"1AF8", x"1C09", x"1CF4", x"1E26", x"1F6F", x"1FC2", x"1F28", x"1E0A", x"1C97", x"1B05", x"19E7", x"18F2", x"17AE", x"160E", x"144E", x"12B2", x"1122", x"0FB5", x"0E8E", x"0DF2", x"0DA4", x"0E09", x"0F19", x"1023", x"1089", x"10B9", x"1038", x"0E57", x"0BAB", x"0964", x"07CC", x"0773", x"0958", x"0C87", x"0F6B", x"11FA", x"148A", x"1626", x"16AC", x"16FB", x"1708", x"1679", x"164C", x"170C", x"179F", x"1790", x"17D5", x"187B", x"18C8", x"191A", x"19C9", x"19CD", x"1935", x"19B5", x"1B2B", x"1C04", x"1C4E", x"1C7B", x"1BAC", x"1A8A", x"1B60", x"1D2E", x"1D6B", x"1CD7", x"1C69", x"1B47", x"1A9F", x"1C8F", x"1EAA", x"1E85", x"1E1B", x"1E32", x"1CBC", x"1AAC", x"1984", x"1747", x"1410", x"1389", x"1588", x"1702", x"1829", x"1976", x"18D7", x"1710", x"16A2", x"1657", x"1472", x"1260", x"111B", x"0FB4", x"0EDB", x"0F7B", x"106C", x"10FD", x"11ED", x"135D", x"145D", x"14B6", x"14CF", x"1521", x"156E", x"15AE", x"15F1", x"156E", x"1372", x"1169", x"10D7", x"10B7", x"1030", x"0FF3", x"0F14", x"0D01", x"0C2C", x"0D93", x"0EFD", x"106C", x"133E", x"15C1", x"16B1", x"1778", x"1759", x"14E2", x"12C2", x"13A5", x"1616", x"198F", x"1E17", x"219D", x"2291", x"22AE", x"226A", x"20C2", x"1E64", x"1C51", x"1A03", x"17CB", x"165C", x"159B", x"1534", x"1534", x"1560", x"15AF", x"15AA", x"14CE", x"141A", x"1454", x"14B6", x"1574", x"171A", x"17BA", x"16CA", x"1697", x"1715", x"162A", x"14D3", x"1389", x"1063", x"0CF4", x"0C80", x"0D3F", x"0CE4", x"0D1E", x"0D9D", x"0C72", x"0B8C", x"0BC2", x"0A02", x"064E", x"03D8", x"02AC", x"0291", x"050E", x"0891", x"0A38", x"0ABF", x"0B1E", x"0A56", x"0985", x"0991", x"091A", x"0798", x"0649", x"04ED", x"03B7", x"0430", x"05C7", x"070E", x"0818", x"08A7", x"0843", x"082F", x"08CF", x"0968", x"0A17", x"0AC5", x"0A0C", x"08BA", x"080A", x"076D", x"072C", x"083F", x"08AC", x"071C", x"05BB", x"04FF", x"03D2", x"03B5", x"051B", x"059B", x"05A2", x"072E", x"0863", x"07FA", x"0787", x"06C3", x"051F", x"0530", x"07E1", x"0B08", x"0EA4", x"12AC", x"14DF", x"1567", x"164C", x"16AC", x"15C7", x"14E3", x"12DC", x"0E71", x"0A70", x"0882", x"0773", x"073F", x"0819", x"0767", x"0501", x"0341", x"0249", x"0197", x"0252", x"0411", x"054A", x"0650", x"0716", x"06CF", x"066F", x"06BB", x"06B8", x"06A7", x"070B", x"06BE", x"060D", x"0663", x"06D2", x"0631", x"063A", x"06C8", x"0637", x"0527", x"0427", x"01AB", x"FEB5", x"FE03", x"FF33", x"0129", x"044E", x"0733", x"07E9", x"0781", x"0719", x"0607", x"04E1", x"0488", x"03B2", x"0219", x"010E", x"0086", x"FFD3", x"FFC2", x"0028", x"FFFA", x"FFCD", x"005A", x"012A", x"01F8", x"0342", x"04CF", x"064B", x"0760", x"0787", x"0698", x"0502", x"0332", x"01F3", x"019E", x"011E", x"FFFE", x"FF27", x"FE5B", x"FCC6", x"FB4E", x"FA96", x"F96C", x"F875", x"F89E", x"F84D", x"F634", x"F439", x"F378", x"F366", x"F54A", x"F939", x"FC73", x"FE06", x"FF84", x"0097", x"00B0", x"00EC", x"00F9", x"FEE4", x"FBD3", x"F9AD", x"F820", x"F74B", x"F83C", x"F933", x"F8B4", x"F7EA", x"F76B", x"F641", x"F551", x"F57B", x"F5A1", x"F5CE", x"F713", x"F82B", x"F7DF", x"F6F7", x"F579", x"F331", x"F1B0", x"F19A", x"F187", x"F18C", x"F1E4", x"F147", x"F023", x"F0A8", x"F24E", x"F3FB", x"F619", x"F73A", x"F581", x"F33E", x"F2EC", x"F3CB", x"F617", x"FA53", x"FDF2", x"FF66", x"00B8", x"01C5", x"0100", x"FFE9", x"FF29", x"FD46", x"FB01", x"FA28", x"F94F", x"F80C", x"F7EE", x"F837", x"F790", x"F749", x"F753", x"F621", x"F4C7", x"F487", x"F46F", x"F4C9", x"F617", x"F66C", x"F491", x"F1B4", x"EE4B", x"EAFD", x"E9AE", x"EA1C", x"EA8B", x"EAD8", x"EA3D", x"E79C", x"E4B5", x"E349", x"E2F3", x"E43D", x"E741", x"E923", x"E8AD", x"E82A", x"E817", x"E868", x"EAF2", x"EF21", x"F225", x"F46B", x"F6F7", x"F832", x"F846", x"F883", x"F7CD", x"F5DC", x"F46B", x"F2F4", x"F0E3", x"EFC9", x"EF5D", x"EE20", x"ED73", x"ED5E", x"EC56", x"EBF7", x"ED71", x"EE18", x"EDF0", x"EF23", x"EFE7", x"EF7C", x"F07C", x"F159", x"EF3D", x"ED39", x"ECDE", x"EBF2", x"EBC0", x"EDAD", x"ED4B", x"EA25", x"E867", x"E7C8", x"E726", x"E990", x"ECE4", x"EBE8", x"E8CA", x"E6E8", x"E4E0", x"E4B7", x"E93D", x"EDC5", x"EF13", x"F02C", x"F0DF", x"EF28", x"EDE6", x"EDB2", x"EB66", x"E831", x"E6CF", x"E55A", x"E3B0", x"E38D", x"E34B", x"E1E5", x"E166", x"E0FC", x"DFD8", x"E021", x"E1B9", x"E2A6", x"E460", x"E6D5", x"E7A6", x"E851", x"EA8F", x"EB4B", x"EA00", x"E940", x"E7A0", x"E4DE", x"E49F", x"E5F7", x"E54B", x"E419", x"E389", x"E188", x"E022", x"E1AD", x"E2D2", x"E219", x"E1D2", x"E146", x"E017", x"E1D4", x"E638", x"EA19", x"EDC0", x"F15E", x"F27C", x"F298", x"F3C9", x"F46D", x"F448", x"F49A", x"F3D0", x"F154", x"EF87", x"EE18", x"EC93", x"ECDF", x"EE37", x"EE4C", x"EEA9", x"EF94", x"EECA", x"EE0C", x"EE9C", x"ED98", x"EBA8", x"EC5F", x"ED95", x"ED79", x"EE69", x"EE50", x"E9FE", x"E60C", x"E557", x"E459", x"E388", x"E4A6", x"E396", x"DFFD", x"DF6E", x"E0E2", x"E0C2", x"E110", x"E1B3", x"DF7A", x"DD75", x"DF16", x"E160", x"E342", x"E6A9", x"E917", x"E91A", x"E9B6", x"EA8F", x"E96C", x"E810", x"E6C8", x"E396", x"E025", x"DE6B", x"DCA7", x"DB58", x"DBF6", x"DC75", x"DC14", x"DCA5", x"DD07", x"DC27", x"DC2A", x"DCEF", x"DCE5", x"DDD2", x"DFD6", x"E050", x"E011", x"DFED", x"DDB1", x"DA3D", x"D908", x"D8ED", x"D8CD", x"DA7D", x"DBAB", x"D94E", x"D697", x"D60A", x"D5B5", x"D647", x"D8B2", x"D968", x"D7AD", x"D7AF", x"D9BD", x"DC5A", x"E096", x"E588", x"E81F", x"E94A", x"EAAD", x"EB4F", x"EB9C", x"ECA2", x"ED04", x"EC2D", x"EB57", x"E9FD", x"E85C", x"E81F", x"E8B5", x"E8E4", x"E979", x"E9EB", x"E91E", x"E89F", x"E927", x"E8F9", x"E8A8", x"E90F", x"E867", x"E70B", x"E716", x"E72C", x"E61B", x"E606", x"E639", x"E518", x"E4E6", x"E639", x"E5BB", x"E3ED", x"E368", x"E2D5", x"E244", x"E467", x"E6E1", x"E5E8", x"E39A", x"E24F", x"E129", x"E22F", x"E6F0", x"EBCC", x"EE5C", x"F027", x"F0DE", x"EF9D", x"EE38", x"ED73", x"EBDD", x"EA26", x"E91F", x"E808", x"E701", x"E6DC", x"E722", x"E7C7", x"E907", x"E9D4", x"EA4D", x"EB3F", x"EC62", x"ED6A", x"EF32", x"F09F", x"F0C6", x"F152", x"F2E7", x"F429", x"F5A9", x"F77B", x"F743", x"F560", x"F45B", x"F3BE", x"F2B1", x"F2FB", x"F417", x"F3E3", x"F3C3", x"F4A4", x"F3B2", x"F0DB", x"EE76", x"ECA7", x"EBAD", x"EE0A", x"F2FA", x"F702", x"F9CE", x"FBCC", x"FBCD", x"FA6D", x"F9B3", x"F943", x"F8A2", x"F8D2", x"F99B", x"F9B9", x"F916", x"F7EE", x"F672", x"F580", x"F5B1", x"F6B8", x"F809", x"F8C5", x"F84A", x"F764", x"F667", x"F522", x"F454", x"F4F3", x"F5F5", x"F73C", x"F94B", x"FA6B", x"F955", x"F7C4", x"F6C5", x"F57D", x"F505", x"F609", x"F687", x"F64C", x"F71E", x"F833", x"F7A2", x"F662", x"F4F9", x"F30A", x"F262", x"F4C5", x"F87D", x"FBD4", x"FEA7", x"0014", x"FF8B", x"FE40", x"FD28", x"FBEE", x"FB0A", x"FABD", x"FA58", x"F967", x"F819", x"F679", x"F538", x"F4F2", x"F5CE", x"F766", x"F918", x"F9BF", x"F945", x"F826", x"F69B", x"F57D", x"F5D4", x"F735", x"F8E1", x"FB48", x"FD42", x"FD1A", x"FB69", x"F95F", x"F6E5", x"F535", x"F5F9", x"F77C", x"F811", x"F8CB", x"FA1C", x"FAB1", x"FAFE", x"FB56", x"FA3B", x"F80D", x"F7B8", x"F9F0", x"FD98", x"0228", x"0691", x"0909", x"09A8", x"099A", x"0948", x"08DE", x"08EF", x"093C", x"095C", x"08F7", x"07F8", x"06E8", x"068C", x"06DB", x"0769", x"07F2", x"0790", x"0610", x"0455", x"02F1", x"01DC", x"017C", x"01DD", x"0265", x"0330", x"04A4", x"0600", x"06C4", x"0709", x"062D", x"042D", x"028A", x"0216", x"0238", x"0316", x"04ED", x"06A5", x"07BA", x"08A5", x"08C2", x"0723", x"04E8", x"040D", x"04D9", x"06EA", x"0A0A", x"0D22", x"0EBC", x"0EF6", x"0EE5", x"0E4D", x"0C9E", x"0AD5", x"09F7", x"095E", x"0891", x"081D", x"077F", x"062C", x"0588", x"067C", x"079D", x"081C", x"08A0", x"08DB", x"08A5", x"0929", x"0A85", x"0B9D", x"0C94", x"0E17", x"0FCC", x"11A0", x"13BC", x"153E", x"153A", x"1423", x"1249", x"105D", x"0F74", x"1047", x"122C", x"14AD", x"16BB", x"1748", x"1616", x"13DC", x"116E", x"1036", x"1101", x"1337", x"164B", x"199D", x"1C2B", x"1DBA", x"1EE1", x"1F21", x"1DEF", x"1C93", x"1BBF", x"1B0C", x"1AEC", x"1B81", x"1B34", x"19B1", x"187A", x"17A6", x"16C3", x"164B", x"166A", x"1609", x"1575", x"155C", x"153A", x"14CF", x"14BC", x"157E", x"16FC", x"18BF", x"1A10", x"1A70", x"1975", x"1724", x"1499", x"12AD", x"1104", x"1070", x"1215", x"14D3", x"16EE", x"182E", x"177F", x"13F4", x"102F", x"0ED8", x"0F93", x"1205", x"168A", x"1AB9", x"1CFC", x"1EBC", x"1FFB", x"1F9B", x"1ED1", x"1E7C", x"1D63", x"1C2A", x"1C02", x"1BB5", x"1AC7", x"1A66", x"19ED", x"18B9", x"186B", x"18DA", x"189B", x"1837", x"17EB", x"1685", x"14FA", x"14CF", x"1519", x"1596", x"173E", x"18B0", x"191E", x"1979", x"194A", x"1777", x"1583", x"13CD", x"119D", x"10BA", x"1283", x"150B", x"1773", x"19AD", x"1909", x"153C", x"11F6", x"10A3", x"10C3", x"139F", x"1897", x"1C4C", x"1EDE", x"219D", x"2326", x"2346", x"23CE", x"2426", x"2395", x"2358", x"2329", x"21DF", x"20A3", x"2016", x"1F54", x"1F1A", x"1FCE", x"1FE3", x"1F84", x"1F68", x"1E6D", x"1C8D", x"1B91", x"1B11", x"1A7D", x"1B18", x"1C83", x"1D4A", x"1E7B", x"2011", x"2074", x"1FF7", x"1F68", x"1DB7", x"1BB8", x"1B81", x"1C37", x"1D9E", x"2097", x"2324", x"22C4", x"2118", x"1F2C", x"1CDD", x"1CD2", x"201C", x"236A", x"255A", x"271A", x"275D", x"263A", x"267C", x"276A", x"26DF", x"25F1", x"24FE", x"2256", x"1FB1", x"1EBF", x"1DBB", x"1C89", x"1C9F", x"1C80", x"1B3D", x"1AB1", x"1A3D", x"1848", x"167E", x"158F", x"1430", x"1372", x"1432", x"1497", x"1493", x"1572", x"15E3", x"158D", x"15D7", x"1599", x"13BD", x"1227", x"1137", x"1008", x"109A", x"133F", x"148B", x"1404", x"12D7", x"102A", x"0D50", x"0DF1", x"1110", x"13CC", x"169C", x"18B8", x"183F", x"1733", x"1763", x"16BD", x"1510", x"140C", x"128A", x"1038", x"0FC6", x"1090", x"1085", x"1099", x"1126", x"1048", x"0ECA", x"0E0D", x"0CC1", x"0AB7", x"09F6", x"0A66", x"0B23", x"0CA6", x"0E38", x"0EF3", x"0F78", x"1026", x"106C", x"10CB", x"1109", x"1041", x"0F5E", x"0EDA", x"0D7C", x"0C4B", x"0D4D", x"0F58", x"10F8", x"12C1", x"1341", x"1125", x"0F50", x"1015", x"11F5", x"145C", x"17A1", x"19A9", x"19BA", x"19C1", x"19DB", x"18EE", x"17EA", x"1721", x"1584", x"1407", x"13B7", x"13C5", x"1400", x"14F4", x"1587", x"14F9", x"145C", x"13A0", x"11F9", x"0FFE", x"0E71", x"0D25", x"0C5D", x"0C7B", x"0D02", x"0DFA", x"0F61", x"1111", x"1307", x"1481", x"1438", x"12C9", x"115F", x"0F0B", x"0C1D", x"0AF2", x"0C02", x"0E0F", x"120B", x"16B4", x"1807", x"15E3", x"13D8", x"12C0", x"124F", x"142D", x"1750", x"18B2", x"1906", x"1A0B", x"1A62", x"199D", x"190E", x"1853", x"16C2", x"15C1", x"157B", x"14F1", x"14B0", x"1513", x"14D8", x"1419", x"1377", x"1221", x"0FE8", x"0E08", x"0C60", x"0A97", x"09E6", x"0A51", x"0ABC", x"0B2E", x"0C00", x"0C93", x"0D02", x"0D5A", x"0CA9", x"0ADA", x"08A0", x"059F", x"0265", x"00BB", x"00A3", x"0168", x"03A9", x"0619", x"05C1", x"0368", x"01ED", x"0109", x"00A7", x"0224", x"03CE", x"0311", x"0192", x"011D", x"002B", x"FE91", x"FE6C", x"FF26", x"FFBA", x"0108", x"02D6", x"02F6", x"01C7", x"00D3", x"001A", x"FF4B", x"FEE5", x"FE6C", x"FD51", x"FC3C", x"FBB3", x"FBB3", x"FC0E", x"FCC9", x"FD94", x"FE7F", x"FFA0", x"0138", x"033B", x"04FB", x"0623", x"06A4", x"062D", x"0498", x"0333", x"02CD", x"034B", x"053F", x"089A", x"0B3E", x"0BAC", x"0B38", x"0A66", x"0948", x"0959", x"0AC3", x"0B98", x"0B8B", x"0BC5", x"0C1F", x"0BF5", x"0C1C", x"0C69", x"0C05", x"0B65", x"0ACC", x"0A04", x"0955", x"0941", x"0998", x"0A5C", x"0B10", x"0AA7", x"0957", x"0813", x"065F", x"04B3", x"0438", x"048A", x"04DF", x"0681", x"08E9", x"0A1B", x"0A4C", x"0A5E", x"090C", x"06D0", x"056C", x"03C2", x"00AE", x"FE5F", x"FDBB", x"FDB9", x"FF8B", x"0325", x"0503", x"03F0", x"0232", x"FFE5", x"FD02", x"FBE9", x"FC7C", x"FC35", x"FBC7", x"FCC5", x"FDAA", x"FDC6", x"FE46", x"FE4F", x"FCDD", x"FB80", x"FAE0", x"F9F3", x"F915", x"F918", x"F916", x"F8D1", x"F899", x"F7CA", x"F5DF", x"F3C1", x"F1A0", x"EF6B", x"EDD0", x"ECE7", x"EBDC", x"EAB6", x"E9BE", x"E8BF", x"E80E", x"E856", x"E90B", x"E943", x"E8AF", x"E70D", x"E465", x"E1B8", x"E005", x"DFA7", x"E0DB", x"E345", x"E5BD", x"E78F", x"E883", x"E878", x"E7D6", x"E742", x"E6FF", x"E6E8", x"E756", x"E852", x"E98A", x"EAA6", x"EBB9", x"EC91", x"ED25", x"ED63", x"ED55", x"ECCC", x"EBC6", x"EABF", x"EA57", x"EA74", x"EAC3", x"EB2B", x"EB70", x"EB3F", x"EAE3", x"EAD8", x"EAA3", x"EA0A", x"E968", x"E8A6", x"E7BB", x"E788", x"E864", x"E998", x"EAF4", x"EC57", x"ECAD", x"EB95", x"EA28", x"E8AD", x"E766", x"E7DF", x"EA8B", x"ED9A", x"F017", x"F20B", x"F265", x"F189", x"F1E3", x"F3C8", x"F5A3", x"F769", x"F970", x"FA55", x"FA86", x"FBB4", x"FCF3", x"FCB2", x"FC50", x"FC5C", x"FBF1", x"FB98", x"FC60", x"FC74", x"FB0E", x"FA13", x"F976", x"F806", x"F660", x"F4DF", x"F232", x"EF1D", x"EDA2", x"ED0E", x"EC85", x"EC7C", x"ECB9", x"EC75", x"EC9B", x"EDAF", x"EE88", x"EECC", x"EE99", x"ED80", x"EBC2", x"EAA5", x"EA4A", x"EAFE", x"ECDE", x"EEC5", x"EF35", x"EEC2", x"EDAA", x"EC3A", x"EBF4", x"ED5C", x"EEA9", x"EF88", x"F09E", x"F10A", x"F088", x"F073", x"F059", x"EF1C", x"EDD1", x"ED46", x"EC09", x"EA83", x"E9C7", x"E915", x"E837", x"E8BD", x"E9F2", x"E9F6", x"E901", x"E777", x"E4B9", x"E217", x"E104", x"E101", x"E113", x"E1BE", x"E2E5", x"E415", x"E578", x"E6E2", x"E787", x"E716", x"E586", x"E358", x"E115", x"DED1", x"DD44", x"DDA1", x"DF62", x"E115", x"E28E", x"E38A", x"E310", x"E264", x"E324", x"E3EA", x"E39A", x"E35E", x"E325", x"E247", x"E270", x"E3FE", x"E4F8", x"E547", x"E5DD", x"E59B", x"E463", x"E3AC", x"E2EE", x"E195", x"E117", x"E15E", x"E127", x"E123", x"E144", x"DFC3", x"DD35", x"DB20", x"D8E5", x"D723", x"D780", x"D8B6", x"D959", x"DAD0", x"DCE4", x"DE74", x"E0B2", x"E3A4", x"E462", x"E2F7", x"E101", x"DE05", x"DB5C", x"DBE0", x"DE48", x"E001", x"E1DF", x"E3AA", x"E3E2", x"E49E", x"E716", x"E897", x"E881", x"E885", x"E805", x"E6D3", x"E73A", x"E8BC", x"E969", x"EA14", x"EB24", x"EB38", x"EB13", x"EBA1", x"EBB5", x"EB81", x"EBE0", x"EBB9", x"EAE5", x"EABE", x"EA8D", x"E97A", x"E8D9", x"E866", x"E72C", x"E700", x"E892", x"E9AC", x"EA69", x"EB85", x"EB76", x"EA77", x"EABA", x"EB06", x"E9A6", x"E7F9", x"E5F5", x"E30D", x"E194", x"E2F1", x"E4E1", x"E6B2", x"E899", x"E8D6", x"E7C9", x"E81B", x"E9A9", x"EB4A", x"EDA1", x"EF9E", x"EF7C", x"EEAE", x"EE23", x"ED03", x"EC42", x"ECC8", x"ECDE", x"ECA6", x"ED8B", x"EE5B", x"EE76", x"EF43", x"EFAE", x"EE1F", x"ECB0", x"EBF5", x"EA5F", x"E921", x"E939", x"E8B8", x"E805", x"E950", x"EB40", x"EC8D", x"EEA6", x"F0C4", x"F14C", x"F220", x"F3B4", x"F3D1", x"F2FE", x"F25E", x"F075", x"EE66", x"EED5", x"F0B3", x"F2B1", x"F592", x"F79A", x"F6DF", x"F5D7", x"F620", x"F66C", x"F77D", x"F9A5", x"F9FE", x"F854", x"F75B", x"F6C5", x"F61C", x"F71E", x"F8E0", x"F92E", x"F952", x"FA23", x"F9EE", x"F96D", x"F9EF", x"FA21", x"FA0A", x"FB46", x"FCD0", x"FD43", x"FD8F", x"FD42", x"FBAC", x"FA5C", x"FA2E", x"FA27", x"FAFD", x"FCBA", x"FDA2", x"FDB5", x"FDA4", x"FC0F", x"F912", x"F66A", x"F318", x"EE8E", x"EBA5", x"EAEF", x"EB17", x"ED62", x"F13F", x"F2B1", x"F197", x"F0FA", x"F0A6", x"F098", x"F2FB", x"F5F0", x"F60C", x"F4FA", x"F4D6", x"F497", x"F4E3", x"F720", x"F8F6", x"F910", x"F93E", x"F9B5", x"F92D", x"F8A6", x"F8BD", x"F859", x"F7E8", x"F80D", x"F7EB", x"F722", x"F62C", x"F50A", x"F423", x"F3E2", x"F3B8", x"F3D7", x"F4BF", x"F583", x"F5A4", x"F608", x"F5CD", x"F451", x"F3B0", x"F43E", x"F3B5", x"F268", x"F1DE", x"F0CB", x"EF7C", x"F08D", x"F264", x"F1F7", x"F0F9", x"F13B", x"F195", x"F300", x"F6F9", x"FA66", x"FAF5", x"FAC5", x"FAC0", x"F9DA", x"F9B6", x"FB93", x"FD8E", x"FF0F", x"0115", x"028D", x"0241", x"0144", x"008D", x"FFE6", x"FFBA", x"FFF7", x"FFF6", x"FF68", x"FEE8", x"FEE2", x"FFDA", x"012B", x"0219", x"02E8", x"03B5", x"0390", x"032A", x"032B", x"026D", x"00E9", x"0074", x"002C", x"FE46", x"FC52", x"FB78", x"FA8B", x"FABB", x"FDB0", x"0066", x"009B", x"00C9", x"0189", x"01B5", x"033B", x"06D2", x"0902", x"0936", x"09FD", x"0AAE", x"09F5", x"09AD", x"09D7", x"0896", x"072B", x"0728", x"06E6", x"05EC", x"056A", x"0502", x"0459", x"0474", x"04C7", x"041F", x"02B3", x"00C2", x"FE58", x"FCB3", x"FC49", x"FC67", x"FD99", x"FF81", x"0077", x"00B4", x"014A", x"0159", x"011A", x"0214", x"028E", x"00FD", x"FF78", x"FEFA", x"FEA1", x"FFEE", x"02FE", x"0440", x"02FB", x"01C8", x"0097", x"FFC3", x"01CA", x"056F", x"076D", x"088E", x"0995", x"0909", x"0830", x"08DE", x"0925", x"0857", x"0872", x"08D8", x"088C", x"095A", x"0AC1", x"0AD4", x"0A91", x"0AF3", x"0AB0", x"0A96", x"0BB7", x"0C2A", x"0BB7", x"0BAE", x"0B4A", x"0A6B", x"0B23", x"0C7D", x"0C85", x"0C8A", x"0C76", x"0AC8", x"09B1", x"0A65", x"09DA", x"0793", x"05C0", x"0346", x"00B5", x"017D", x"0451", x"0587", x"062C", x"06D7", x"05E8", x"05C6", x"08AC", x"0B8A", x"0CE4", x"0E57", x"0E36", x"0BFF", x"0B3D", x"0C33", x"0C5E", x"0D50", x"0F53", x"0FC9", x"0FAD", x"1134", x"120B", x"116E", x"11DB", x"1274", x"1217", x"12B6", x"141C", x"13EA", x"1338", x"1312", x"121F", x"1153", x"11ED", x"127E", x"12FF", x"1466", x"1514", x"1490", x"14F3", x"154B", x"146D", x"13F3", x"1375", x"112A", x"0FAA", x"1097", x"114B", x"1191", x"1289", x"1223", x"1074", x"112C", x"13B6", x"15CD", x"187A", x"1AB7", x"19C5", x"1786", x"163E", x"1476", x"1325", x"1418", x"151B", x"1517", x"162B", x"177A", x"172F", x"173A", x"1799", x"1683", x"157E", x"15DC", x"15A2", x"155E", x"1652", x"16D2", x"1696", x"1787", x"184F", x"17F5", x"1887", x"18F1", x"171D", x"157F", x"151A", x"13A9", x"1270", x"12E4", x"11F2", x"0FBB", x"1003", x"11BD", x"1262", x"13AB", x"14CC", x"133E", x"11E3", x"13A2", x"15EA", x"17CB", x"1A2C", x"1A7F", x"17D4", x"156C", x"13CB", x"11A3", x"1089", x"10E7", x"10A7", x"10A5", x"1224", x"1360", x"13D0", x"1483", x"149C", x"13D7", x"13D3", x"145B", x"1480", x"14FB", x"158D", x"154F", x"154F", x"15CB", x"15E3", x"1693", x"1862", x"1979", x"19CE", x"1A9D", x"1AD3", x"1A57", x"1AEE", x"1BC1", x"1B31", x"1AC9", x"1B89", x"1BF0", x"1C5E", x"1D29", x"1CBB", x"1B2C", x"1A9D", x"1B1A", x"1C41", x"1E8F", x"20E6", x"21CF", x"2202", x"21AA", x"2061", x"1FB8", x"2053", x"20DD", x"2160", x"2255", x"2293", x"2235", x"22BE", x"2341", x"22B6", x"2254", x"2216", x"214B", x"216B", x"22DB", x"23B3", x"2419", x"24D8", x"24C8", x"244B", x"2561", x"26C6", x"2677", x"2593", x"243A", x"2157", x"1EF5", x"1E84", x"1DC2", x"1BD8", x"1A80", x"1996", x"184D", x"1826", x"18B3", x"17F8", x"1685", x"15FB", x"15F4", x"1663", x"17B7", x"18F3", x"18EE", x"1842", x"16E7", x"14DA", x"1314", x"123A", x"11D8", x"11D9", x"124A", x"124F", x"11DA", x"1181", x"1103", x"1027", x"0F69", x"0F12", x"0EC4", x"0EB0", x"0ED5", x"0EF5", x"0EF3", x"0F02", x"0EF6", x"0ED0", x"0EAC", x"0E7E", x"0E54", x"0E50", x"0E4C", x"0E29", x"0E11", x"0DF9", x"0D7D", x"0C8B", x"0B8D", x"0AAD", x"09D9", x"0921", x"08AA", x"085B", x"085C", x"095D", x"0B69", x"0DC7", x"1002", x"123F", x"13F0", x"1477", x"13F3", x"12B0", x"10BF", x"0EDA", x"0DFE", x"0DD6", x"0D7B", x"0CE5", x"0C58", x"0BAD", x"0B37", x"0B7F", x"0BF9", x"0C3B", x"0CBD", x"0DCC", x"0F0F", x"1085", x"123C", x"1358", x"137D", x"1351", x"1300", x"1237", x"117D", x"113C", x"10F3", x"10AD", x"1134", x"11FE", x"1235", x"127E", x"136B", x"1479", x"15BC", x"1770", x"187E", x"183F", x"181A", x"18BC", x"19CF", x"1B4F", x"1CF9", x"1D79", x"1CA3", x"1B5E", x"19A3", x"176C", x"1574", x"13C3", x"121B", x"1134", x"114B", x"11B6", x"1260", x"133E", x"134D", x"1295", x"11F7", x"1165", x"10EF", x"1132", x"11A7", x"1155", x"10BA", x"0FF3", x"0EAC", x"0D84", x"0D1C", x"0C93", x"0BD4", x"0BC4", x"0BE9", x"0BD7", x"0C72", x"0D1E", x"0CB4", x"0BD9", x"0B89", x"0AE7", x"09F4", x"095C", x"085A", x"06A6", x"05E0", x"06A3", x"07EF", x"09A4", x"0B84", x"0C73", x"0C2F", x"0B5E", x"09D5", x"0782", x"052A", x"0339", x"01D5", x"0148", x"0167", x"01C3", x"023C", x"029A", x"0281", x"022E", x"01C3", x"014C", x"014F", x"01EE", x"02A4", x"0323", x"034F", x"0295", x"018C", x"0113", x"011B", x"0118", x"0150", x"012A", x"000D", x"FF37", x"FF44", x"FF3F", x"FEE8", x"FED6", x"FE53", x"FD2E", x"FC7B", x"FC0C", x"FACF", x"F986", x"F919", x"F948", x"FA38", x"FC2A", x"FE41", x"FF8B", x"0042", x"0010", x"FED4", x"FD43", x"FBCA", x"FAA3", x"FA2F", x"FA3C", x"FA25", x"FA00", x"FA14", x"F9CF", x"F973", x"F96F", x"F942", x"F8D5", x"F8E6", x"F90C", x"F8D6", x"F8D2", x"F906", x"F8EA", x"F8F2", x"F988", x"F9A5", x"F959", x"F920", x"F888", x"F760", x"F6D7", x"F6B9", x"F5FC", x"F535", x"F4D4", x"F42E", x"F356", x"F33B", x"F2DA", x"F1D4", x"F173", x"F28D", x"F49B", x"F787", x"FAF5", x"FD71", x"FE7E", x"FEB0", x"FE3D", x"FD04", x"FB5C", x"F9AF", x"F7F9", x"F686", x"F54D", x"F44D", x"F375", x"F2C8", x"F24B", x"F236", x"F24D", x"F239", x"F252", x"F2AE", x"F321", x"F3B2", x"F499", x"F534", x"F54D", x"F56F", x"F57B", x"F4FB", x"F442", x"F39F", x"F268", x"F11B", x"F089", x"F03D", x"EFA7", x"EF74", x"EFC6", x"EFF1", x"F042", x"F0F5", x"F123", x"F0A6", x"F0DE", x"F25C", x"F473", x"F6EB", x"F91F", x"F9EA", x"F8F7", x"F795", x"F619", x"F47E", x"F302", x"F1E2", x"F0AA", x"EF4F", x"EE3B", x"ED92", x"ED25", x"ED1E", x"ED76", x"ED95", x"ED2A", x"EC3E", x"EB70", x"EAF7", x"EB26", x"EBF9", x"ECDD", x"ECFE", x"EC6F", x"EBCC", x"EB1F", x"EA75", x"EA2D", x"E9E9", x"E941", x"E8EB", x"E996", x"EAAB", x"EBB4", x"ED09", x"EE39", x"EE83", x"EE66", x"EE44", x"ED4A", x"EC15", x"EC3A", x"EDD5", x"F012", x"F2D3", x"F576", x"F6D2", x"F732", x"F793", x"F7AF", x"F725", x"F65D", x"F58D", x"F499", x"F40C", x"F42C", x"F4DF", x"F5CB", x"F6E5", x"F7B7", x"F837", x"F819", x"F79F", x"F75C", x"F792", x"F7F4", x"F88C", x"F940", x"F941", x"F8CA", x"F88D", x"F7F5", x"F68B", x"F4F4", x"F330", x"F0C9", x"EF13", x"EED3", x"EED0", x"EEDA", x"EFEF", x"F13E", x"F1B6", x"F23B", x"F25E", x"F0B4", x"EE9A", x"EE13", x"EE7F", x"EF45", x"F0E8", x"F234", x"F1F7", x"F199", x"F1D5", x"F1C2", x"F145", x"F0E9", x"F029", x"EEF7", x"EE59", x"EE47", x"EE3D", x"EE82", x"EED6", x"EED0", x"EEB1", x"EE84", x"EE31", x"EE12", x"EE36", x"EE3F", x"EE66", x"EEEE", x"EF45", x"EFAE", x"F074", x"F0C0", x"F047", x"EFCF", x"EF0B", x"EDD0", x"ED43", x"ED58", x"ECD9", x"EC3E", x"EC4A", x"EC1A", x"EB84", x"EB70", x"EAE5", x"E91B", x"E7C9", x"E807", x"E91A", x"EB1B", x"EE04", x"F030", x"F0DF", x"F109", x"F0C1", x"EFDB", x"EF12", x"EE83", x"EDBF", x"EC96", x"EB30", x"E990", x"E86F", x"E849", x"E8C1", x"E9EE", x"EB56", x"EC3B", x"ECF1", x"EE14", x"EEEB", x"EF5A", x"EFE2", x"EFFE", x"EF20", x"EE73", x"EDC7", x"EC46", x"EA8E", x"E961", x"E7CA", x"E675", x"E6AB", x"E772", x"E7EB", x"E948", x"EB38", x"EC67", x"EDA4", x"EF33", x"EF24", x"EDD4", x"ED7B", x"EE0E", x"EF21", x"F17F", x"F412", x"F49F", x"F3CE", x"F2D7", x"F164", x"EFE1", x"EF2F", x"EE65", x"ECC1", x"EB12", x"E979", x"E7D0", x"E6F3", x"E6E8", x"E6BE", x"E672", x"E632", x"E593", x"E50B", x"E549", x"E5C9", x"E64F", x"E75C", x"E866", x"E8DD", x"E90C", x"E8D0", x"E77C", x"E5F5", x"E47A", x"E2CA", x"E145", x"E0A5", x"E036", x"E010", x"E0DB", x"E1E3", x"E24E", x"E293", x"E24D", x"E0A9", x"DEFB", x"DEDA", x"E012", x"E2A1", x"E679", x"E9E9", x"EB81", x"EC10", x"EC29", x"EB89", x"EADC", x"EA83", x"E9B1", x"E864", x"E759", x"E6A4", x"E660", x"E721", x"E8A2", x"EA35", x"EBA3", x"ECB2", x"ED09", x"ED2C", x"ED56", x"ED53", x"ED45", x"ED20", x"EC92", x"EBCF", x"EB54", x"EAC8", x"EA19", x"E99F", x"E888", x"E6E2", x"E59F", x"E506", x"E483", x"E4CA", x"E5E6", x"E686", x"E6F0", x"E7E0", x"E80A", x"E6DE", x"E60C", x"E603", x"E664", x"E841", x"EBAA", x"EE28", x"EF4E", x"F066", x"F100", x"F0D6", x"F140", x"F1BB", x"F0D6", x"EF4B", x"EE1E", x"EC7B", x"EB07", x"EAB5", x"EAC3", x"EAB0", x"EB59", x"EC7C", x"ED51", x"EE80", x"F012", x"F0FE", x"F1D6", x"F31C", x"F435", x"F533", x"F6A0", x"F77A", x"F75A", x"F70D", x"F625", x"F467", x"F2D2", x"F179", x"EFB1", x"EE68", x"EE3F", x"EE0D", x"EDE1", x"EE1F", x"ED75", x"EBC1", x"EB17", x"EBC2", x"ED49", x"F037", x"F3D6", x"F59D", x"F5E4", x"F5EA", x"F571", x"F49A", x"F4BA", x"F4D3", x"F3BC", x"F2B4", x"F211", x"F123", x"F07A", x"F0A4", x"F0A0", x"F069", x"F0D7", x"F14A", x"F166", x"F1BD", x"F1FA", x"F1B0", x"F178", x"F13C", x"F095", x"F028", x"EFEC", x"EF3A", x"EE89", x"EE45", x"EDA3", x"ED1A", x"ED79", x"ED9E", x"ED48", x"EDA1", x"EE51", x"EE6E", x"EEEE", x"EF7D", x"EE9A", x"ED49", x"ED2E", x"EDDD", x"EF97", x"F2E2", x"F5C4", x"F669", x"F5E7", x"F495", x"F28A", x"F1AB", x"F25D", x"F2CD", x"F2AE", x"F291", x"F18F", x"F026", x"F000", x"F065", x"F03D", x"F080", x"F0F6", x"F0CE", x"F0FF", x"F216", x"F2C2", x"F355", x"F496", x"F59A", x"F675", x"F810", x"F96D", x"F9D0", x"FA34", x"FA42", x"F953", x"F903", x"F9BA", x"F9FA", x"FA50", x"FBB7", x"FCA7", x"FD0D", x"FE55", x"FF06", x"FDED", x"FD04", x"FD32", x"FDCB", x"FFE9", x"03C9", x"06AB", x"07ED", x"08DA", x"0909", x"08B6", x"09A0", x"0B3E", x"0BDE", x"0C67", x"0D09", x"0CFC", x"0D68", x"0F2E", x"10C6", x"1189", x"1269", x"128D", x"11B3", x"1146", x"111A", x"1037", x"0F84", x"0F69", x"0F13", x"0F09", x"0FBE", x"0FF3", x"0FAC", x"0F73", x"0EAB", x"0D4A", x"0CE0", x"0CE5", x"0CAE", x"0CFF", x"0DB1", x"0D6C", x"0D0B", x"0D0B", x"0BDA", x"09AB", x"082E", x"0747", x"06E4", x"0843", x"0A45", x"0ADE", x"0A5F", x"096F", x"07B0", x"0641", x"0664", x"06CC", x"06A6", x"066B", x"058E", x"03F1", x"02E3", x"02AE", x"024A", x"0203", x"01FC", x"017D", x"0104", x"013A", x"01B0", x"0256", x"0382", x"0473", x"04D9", x"0581", x"0603", x"0626", x"0680", x"0695", x"055D", x"040E", x"036E", x"0270", x"016B", x"0151", x"0116", x"0082", x"0126", x"025D", x"025C", x"020C", x"0255", x"0284", x"0378", x"0645", x"08F1", x"0A08", x"0A1E", x"0911", x"06B4", x"0504", x"04AE", x"0468", x"041C", x"0404", x"033F", x"0210", x"01ED", x"025D", x"02B0", x"039A", x"04DE", x"0599", x"066A", x"077B", x"082D", x"08C1", x"099D", x"09FA", x"09E1", x"09DF", x"098D", x"08D7", x"0876", x"07CF", x"0685", x"05E0", x"064A", x"06A0", x"077D", x"0959", x"0AED", x"0C02", x"0DB4", x"0EE1", x"0E76", x"0DED", x"0E74", x"0FA1", x"11E1", x"157C", x"1852", x"1945", x"18F7", x"17CC", x"15EB", x"148F", x"1425", x"1416", x"1442", x"1483", x"147C", x"1448", x"1456", x"1463", x"1491", x"14E7", x"150C", x"150D", x"1585", x"1651", x"1760", x"18EC", x"1A50", x"1AFC", x"1B66", x"1BBA", x"1B71", x"1B10", x"1AA5", x"1930", x"170D", x"1580", x"145B", x"1364", x"139F", x"14AA", x"1542", x"15CD", x"1694", x"1637", x"14DA", x"13FD", x"1410", x"1506", x"177D", x"1A81", x"1C5B", x"1CAB", x"1BCB", x"19DF", x"17DD", x"169B", x"15D5", x"1578", x"155B", x"1492", x"1344", x"1293", x"1283", x"12C2", x"13D8", x"1521", x"155F", x"1558", x"15D9", x"15ED", x"1596", x"15CA", x"15DF", x"1579", x"15D1", x"16AA", x"16A3", x"1621", x"15BC", x"1479", x"12EC", x"126C", x"123E", x"1190", x"117F", x"11F3", x"11CB", x"117C", x"116D", x"1027", x"0DE5", x"0C92", x"0CA5", x"0DC0", x"1019", x"131F", x"1531", x"162C", x"16C4", x"16D8", x"1672", x"163A", x"1640", x"165C", x"1631", x"1557", x"13BD", x"11F3", x"1052", x"0EFF", x"0E56", x"0E1B", x"0DE4", x"0E27", x"0F1B", x"1007", x"10D0", x"11EB", x"1353", x"14C7", x"16B1", x"18A7", x"19E2", x"1A5A", x"1A3F", x"195B", x"17F5", x"16B8", x"1583", x"145B", x"13B3", x"1366", x"1315", x"12E0", x"12B8", x"1207", x"1143", x"1187", x"1302", x"155C", x"1861", x"1B1A", x"1C96", x"1CAE", x"1BD2", x"1A49", x"186F", x"16CA", x"15B3", x"14F4", x"1406", x"129E", x"1142", x"103F", x"0F7D", x"0F3B", x"0F6B", x"0F48", x"0EE1", x"0F30", x"0FF8", x"107A", x"10F4", x"1195", x"11A2", x"1193", x"1218", x"1295", x"127F", x"1296", x"128E", x"11F3", x"1177", x"116B", x"10E0", x"103B", x"102F", x"0FFE", x"0F66", x"0F01", x"0DFC", x"0BAD", x"0996", x"0935", x"0A35", x"0CEA", x"1122", x"14A1", x"163E", x"16AE", x"1666", x"1563", x"14E8", x"1546", x"15BF", x"1624", x"166B", x"15FB", x"14CA", x"1378", x"11B8", x"0FC1", x"0E16", x"0CA1", x"0B47", x"0AB3", x"0A9C", x"0A29", x"09CA", x"09D8", x"09D6", x"0A1B", x"0B32", x"0C31", x"0CAA", x"0D10", x"0D33", x"0C89", x"0BE8", x"0B82", x"0AEB", x"0AA9", x"0B39", x"0BC2", x"0C05", x"0C20", x"0B85", x"0A08", x"091A", x"0979", x"0AD5", x"0D28", x"0FE1", x"11A4", x"1212", x"11BF", x"10FB", x"1003", x"0F52", x"0F42", x"0FE2", x"1102", x"124B", x"13B1", x"1512", x"1614", x"16D0", x"179F", x"17EC", x"1778", x"1740", x"174E", x"16E3", x"1645", x"15C2", x"147C", x"1319", x"130C", x"13E2", x"14BA", x"15E0", x"168B", x"15AF", x"1462", x"13D2", x"134A", x"12E1", x"1359", x"1394", x"12C6", x"11F1", x"10D7", x"0E67", x"0BBD", x"0A3F", x"09C8", x"0AAA", x"0D6F", x"1086", x"1244", x"12F4", x"12C4", x"119E", x"1073", x"1007", x"0FFB", x"102C", x"1093", x"1091", x"0FDB", x"0EA9", x"0CE0", x"0AC1", x"08D7", x"0722", x"05A4", x"04F5", x"04F0", x"04F3", x"052B", x"0596", x"05D0", x"0614", x"0703", x"0804", x"0899", x"0903", x"092E", x"089B", x"07E0", x"0729", x"062B", x"04F8", x"0454", x"043D", x"0424", x"0433", x"042D", x"039A", x"02EB", x"0343", x"04AD", x"0672", x"0855", x"09DD", x"0A18", x"090A", x"07AE", x"0602", x"03BE", x"01EC", x"0172", x"01A9", x"0251", x"038E", x"0457", x"03EF", x"038A", x"03F1", x"046B", x"04F2", x"05E5", x"067A", x"0641", x"0621", x"061A", x"057D", x"04C2", x"0472", x"042D", x"03F7", x"041A", x"0418", x"0365", x"0248", x"010F", x"FFD8", x"FF2B", x"FF30", x"FFB4", x"003D", x"006D", x"FFEA", x"FEDE", x"FDA1", x"FCCD", x"FD27", x"FEC9", x"0125", x"03C3", x"0605", x"071F", x"071D", x"0676", x"0528", x"0376", x"022E", x"015E", x"00BF", x"00A0", x"00CA", x"005B", x"FF63", x"FE08", x"FC07", x"F9E3", x"F866", x"F789", x"F727", x"F77B", x"F806", x"F857", x"F8AE", x"F8FD", x"F8D3", x"F8CB", x"F8EF", x"F8C6", x"F87D", x"F85C", x"F764", x"F5E4", x"F4A8", x"F379", x"F25C", x"F289", x"F336", x"F2F1", x"F224", x"F119", x"EF4F", x"EE3E", x"EF5E", x"F14A", x"F305", x"F518", x"F680", x"F661", x"F62B", x"F63C", x"F518", x"F3D1", x"F361", x"F2FA", x"F2E6", x"F473", x"F629", x"F6AB", x"F702", x"F701", x"F5EA", x"F55E", x"F612", x"F64B", x"F60A", x"F62F", x"F5B9", x"F492", x"F434", x"F435", x"F39E", x"F37A", x"F3E4", x"F3C3", x"F357", x"F306", x"F1BD", x"EFE2", x"EEA5", x"EDBC", x"ED21", x"ED67", x"ED8C", x"ECAC", x"EB5B", x"E9F4", x"E84C", x"E7DD", x"E90C", x"EAC6", x"ED02", x"EFB5", x"F18E", x"F289", x"F36C", x"F37A", x"F24A", x"F11D", x"EFB6", x"EDCC", x"ECCD", x"ECFE", x"ECA7", x"EBDA", x"EAD0", x"E895", x"E5CF", x"E4AF", x"E4E6", x"E571", x"E6DE", x"E887", x"E934", x"E9DB", x"EB44", x"ECAB", x"EE2C", x"F044", x"F1B8", x"F24A", x"F295", x"F1F7", x"F06A", x"EF0E", x"ED98", x"EB94", x"EA52", x"E9D3", x"E8B9", x"E782", x"E6B8", x"E52D", x"E3D5", x"E4C5", x"E706", x"E95D", x"EC66", x"EF15", x"F000", x"F096", x"F1BB", x"F1D9", x"F139", x"F0FC", x"EFEF", x"EE5C", x"EE3D", x"EEE4", x"EED3", x"EEC2", x"EE8D", x"ECF1", x"EB5A", x"EB45", x"EB4B", x"EAF7", x"EB10", x"EAE3", x"E9E0", x"E966", x"E990", x"E971", x"E994", x"EA27", x"EA83", x"EAC7", x"EB25", x"EAF1", x"EA97", x"EA9B", x"EA3F", x"E9AF", x"E9C8", x"E9B1", x"E8C0", x"E7EA", x"E699", x"E42C", x"E26A", x"E2A8", x"E3A9", x"E528", x"E77B", x"E8FD", x"E929", x"E999", x"EA13", x"E980", x"E8A2", x"E7FD", x"E6E0", x"E64B", x"E70B", x"E7E9", x"E838", x"E846", x"E753", x"E528", x"E366", x"E264", x"E1D3", x"E22C", x"E325", x"E38A", x"E398", x"E40A", x"E469", x"E50D", x"E676", x"E7B4", x"E849", x"E8E4", x"E92D", x"E8EB", x"E922", x"E9AF", x"E951", x"E8D0", x"E89F", x"E7FB", x"E716", x"E6EC", x"E687", x"E5A6", x"E5F9", x"E779", x"E90B", x"EAE7", x"ECF8", x"EE2A", x"EEEB", x"F04E", x"F15F", x"F1B2", x"F1D6", x"F1AC", x"F115", x"F16F", x"F2E2", x"F478", x"F609", x"F744", x"F70A", x"F5D7", x"F509", x"F490", x"F438", x"F449", x"F41D", x"F2F2", x"F1A8", x"F0D0", x"F05C", x"F09A", x"F1D3", x"F326", x"F43C", x"F515", x"F549", x"F4FB", x"F4E5", x"F4E3", x"F4C8", x"F4ED", x"F502", x"F468", x"F351", x"F1F6", x"EFF3", x"EE01", x"ECE0", x"EC6E", x"EC7C", x"ED69", x"EEA2", x"EFB3", x"F0A4", x"F141", x"F104", x"F062", x"EFAD", x"EEAC", x"EDE2", x"EDDF", x"EE2E", x"EE85", x"EED9", x"EE85", x"ED05", x"EB48", x"EA01", x"E92C", x"E8EB", x"E96E", x"E9ED", x"EA22", x"EA7B", x"EAE7", x"EB6A", x"EC09", x"ECC2", x"ED5D", x"EDA6", x"ED92", x"ED18", x"EC89", x"EC01", x"EB70", x"EB2A", x"EADE", x"EA4F", x"E9A7", x"E955", x"E931", x"E944", x"E9EF", x"EADB", x"EBCB", x"ECF2", x"EE3A", x"EF10", x"EF84", x"EFB7", x"EF72", x"EEC5", x"EE33", x"EDAB", x"ED18", x"ECF8", x"ED59", x"EDC0", x"EE21", x"EE65", x"EE2F", x"ED75", x"ECE8", x"ECD3", x"ED17", x"ED86", x"EE25", x"EE61", x"EE0E", x"ED97", x"ED61", x"ED3A", x"ED5E", x"EE20", x"EF33", x"EFD0", x"F003", x"EFE6", x"EF77", x"EF22", x"EFAB", x"F099", x"F0F1", x"F0D3", x"F04F", x"EF63", x"EE9C", x"EEA3", x"EF1F", x"EFA4", x"F058", x"F120", x"F1A8", x"F248", x"F32E", x"F423", x"F4DF", x"F55B", x"F542", x"F4AD", x"F401", x"F3BA", x"F428", x"F524", x"F632", x"F6DE", x"F6E5", x"F634", x"F543", x"F4AE", x"F47D", x"F492", x"F525", x"F5DF", x"F62E", x"F653", x"F67B", x"F632", x"F5DC", x"F5E7", x"F5B5", x"F4F1", x"F422", x"F36A", x"F2BD", x"F2F8", x"F436", x"F579", x"F63D", x"F688", x"F607", x"F520", x"F4F8", x"F5A0", x"F6D2", x"F879", x"FA0B", x"FB12", x"FBD9", x"FC7F", x"FCE3", x"FD79", x"FE16", x"FDF8", x"FD70", x"FD1E", x"FCC0", x"FCD2", x"FDFE", x"FEFA", x"FECC", x"FE5C", x"FDE1", x"FCDF", x"FC70", x"FD0C", x"FD42", x"FD37", x"FDF7", x"FEBC", x"FEE2", x"FF6C", x"000F", x"FFCD", x"FFD3", x"0074", x"00B1", x"008A", x"00B4", x"0022", x"FEE6", x"FE3C", x"FDCB", x"FCB8", x"FBB3", x"FA9C", x"F8A8", x"F70D", x"F692", x"F69B", x"F6F7", x"F821", x"F903", x"F989", x"FA75", x"FBCE", x"FD2C", x"FF23", x"00F0", x"0185", x"0154", x"00BC", x"FF81", x"FEB9", x"FEDB", x"FE93", x"FDAC", x"FCD1", x"FB92", x"F9F1", x"F94B", x"F94A", x"F8E4", x"F8BF", x"F901", x"F8D7", x"F8E2", x"F9E1", x"FAD4", x"FBB0", x"FD33", x"FE96", x"FF51", x"009B", x"01DF", x"0258", x"02FB", x"043E", x"04D4", x"0515", x"0595", x"050D", x"0394", x"02BE", x"0288", x"0265", x"031E", x"0440", x"04A6", x"04D4", x"0530", x"053D", x"0583", x"0689", x"0746", x"0786", x"07D7", x"07AA", x"070F", x"0777", x"0848", x"0840", x"07F7", x"07B9", x"06BD", x"0612", x"06B3", x"073F", x"073C", x"0794", x"07E4", x"079B", x"07DB", x"0893", x"08AA", x"08C0", x"095C", x"09A5", x"09BC", x"0A43", x"0A67", x"09E3", x"09CB", x"09F5", x"09AF", x"095F", x"08C8", x"0742", x"059D", x"04F0", x"0515", x"060E", x"07DA", x"095B", x"0A0C", x"0A57", x"0A66", x"0A72", x"0B51", x"0CAE", x"0D7E", x"0DC9", x"0D79", x"0C5F", x"0B7C", x"0BB1", x"0C2F", x"0C79", x"0CC3", x"0C74", x"0B4A", x"0A59", x"09BD", x"08DD", x"0818", x"07A6", x"06F6", x"0638", x"062A", x"063F", x"061D", x"065B", x"06B5", x"06B9", x"06EE", x"07A5", x"0825", x"08A9", x"09E0", x"0B47", x"0C1D", x"0C76", x"0C28", x"0AD5", x"0973", x"0933", x"09E5", x"0AD5", x"0BDF", x"0CCE", x"0D47", x"0D94", x"0E17", x"0EB1", x"0EEE", x"0F04", x"0F4C", x"0F85", x"0F7B", x"0F89", x"1010", x"10FA", x"1227", x"137F", x"1475", x"14A7", x"1476", x"148D", x"14E1", x"154D", x"15E1", x"1672", x"16BA", x"16E5", x"1741", x"1787", x"179E", x"1799", x"1758", x"16B4", x"161A", x"15C8", x"1555", x"14EC", x"14C2", x"1480", x"13CE", x"12F5", x"11E8", x"106B", x"0F97", x"1039", x"11AD", x"1350", x"150E", x"165F", x"16F4", x"17A8", x"18C2", x"19AB", x"1A54", x"1AF9", x"1B1E", x"1ABF", x"1A2C", x"1973", x"18BF", x"185A", x"17FB", x"173D", x"1680", x"15B5", x"14C5", x"1439", x"141A", x"13B7", x"136E", x"13BF", x"1415", x"1465", x"1553", x"1684", x"177B", x"18EA", x"1AA4", x"1B8B", x"1BF6", x"1C5F", x"1C48", x"1C1D", x"1CBC", x"1D39", x"1C8A", x"1B24", x"1934", x"16B5", x"1501", x"14D1", x"151B", x"156A", x"15CA", x"15AE", x"1519", x"14F7", x"1525", x"156B", x"1618", x"16C8", x"16FF", x"1741", x"17E1", x"1852", x"1907", x"1A02", x"1A3C", x"19B4", x"1958", x"18E5", x"1838", x"182C", x"186D", x"1827", x"17F4", x"1813", x"17AB", x"16FE", x"16C4", x"162F", x"1571", x"1582", x"15E7", x"15EC", x"164A", x"16D2", x"1683", x"1613", x"1637", x"15DD", x"14E7", x"1449", x"13CE", x"132F", x"139F", x"1531", x"16A8", x"17EA", x"1939", x"19F5", x"1A15", x"1A3A", x"1A56", x"1A64", x"1AD5", x"1B85", x"1BE5", x"1BC8", x"1B1C", x"1A00", x"190A", x"1862", x"17AC", x"1705", x"167D", x"15C4", x"151C", x"14C9", x"1448", x"1394", x"1318", x"12B2", x"1212", x"11CD", x"1203", x"1234", x"12B2", x"137D", x"13DB", x"13A7", x"1374", x"1346", x"1307", x"1366", x"1420", x"141E", x"1336", x"11B0", x"0F97", x"0DBE", x"0D13", x"0D6F", x"0E10", x"0EC0", x"0F67", x"0FBD", x"101C", x"10C9", x"119A", x"1284", x"1371", x"142D", x"14AD", x"1514", x"1578", x"160F", x"16EE", x"1775", x"1755", x"16BF", x"15BD", x"145A", x"131E", x"1258", x"1196", x"111B", x"1140", x"1195", x"11B1", x"11D2", x"11C7", x"1150", x"111A", x"1188", x"121A", x"12C4", x"1379", x"13A7", x"1338", x"1323", x"1308", x"1258", x"1168", x"1064", x"0EFB", x"0DF7", x"0E4D", x"0F13", x"0F60", x"0FB6", x"0FF0", x"0F77", x"0EFC", x"0F11", x"0EEA", x"0E88", x"0EB8", x"0F2E", x"0F1E", x"0EA8", x"0DF6", x"0CC5", x"0BDF", x"0BCB", x"0C1F", x"0C5C", x"0C4D", x"0BAE", x"0A9A", x"0986", x"0892", x"07A2", x"070D", x"06A8", x"0653", x"0657", x"06B1", x"071A", x"07BB", x"0875", x"08A6", x"0870", x"0845", x"080C", x"07F2", x"0884", x"0917", x"08D6", x"082B", x"076F", x"0639", x"056C", x"0594", x"05DD", x"05CE", x"0613", x"0656", x"0633", x"0635", x"0694", x"0679", x"0634", x"0640", x"060D", x"05A1", x"0587", x"05AB", x"05C6", x"0664", x"0727", x"0771", x"0772", x"0755", x"06BD", x"0610", x"05CA", x"058B", x"0568", x"05A6", x"05B5", x"053C", x"04AE", x"0411", x"0330", x"02B4", x"029D", x"0233", x"01CD", x"01CE", x"01BB", x"019A", x"01C0", x"018F", x"0097", x"FFD4", x"FFA1", x"FFE5", x"0123", x"0300", x"0428", x"045C", x"03FE", x"02CA", x"014B", x"008A", x"0006", x"FF33", x"FEBC", x"FE79", x"FDB9", x"FD1E", x"FD13", x"FC86", x"FBA7", x"FB73", x"FB6D", x"FB37", x"FB68", x"FBCC", x"FB78", x"FB10", x"FB12", x"FABB", x"FA2E", x"F9DE", x"F942", x"F88E", x"F891", x"F8E4", x"F90E", x"F96F", x"F9A5", x"F917", x"F881", x"F863", x"F81F", x"F7F5", x"F862", x"F86E", x"F7D9", x"F797", x"F7BD", x"F7E1", x"F8CC", x"FA61", x"FB8F", x"FC80", x"FDC4", x"FEAE", x"FF1F", x"FFEB", x"00A9", x"0108", x"019C", x"0256", x"0281", x"025D", x"0264", x"024D", x"021B", x"021F", x"01DC", x"0148", x"00C3", x"0051", x"FFE7", x"FFCC", x"FFB2", x"FF8C", x"FFCD", x"0041", x"005F", x"008A", x"00C1", x"007E", x"0050", x"00B0", x"00D3", x"007C", x"006C", x"002D", x"FF67", x"FEDB", x"FE46", x"FC9E", x"FA96", x"F931", x"F835", x"F80A", x"F956", x"FAAE", x"FB08", x"FB14", x"FAF3", x"FA44", x"FA15", x"FAC1", x"FB1E", x"FB50", x"FBD5", x"FBF5", x"FB76", x"FB3E", x"FADE", x"F9E2", x"F92A", x"F8B0", x"F7C3", x"F6E8", x"F67C", x"F596", x"F463", x"F3A0", x"F2B9", x"F19B", x"F12C", x"F10D", x"F095", x"F085", x"F0F9", x"F129", x"F1B1", x"F2C2", x"F346", x"F356", x"F3CF", x"F40F", x"F3DA", x"F3EE", x"F3B5", x"F269", x"F140", x"F10B", x"F103", x"F169", x"F26A", x"F2C1", x"F241", x"F228", x"F252", x"F262", x"F2EB", x"F383", x"F32C", x"F293", x"F21A", x"F152", x"F0C0", x"F10D", x"F140", x"F0FA", x"F109", x"F0F4", x"F07F", x"F09C", x"F146", x"F172", x"F162", x"F182", x"F131", x"F0AF", x"F0A1", x"F054", x"EF98", x"EF08", x"EE6A", x"EDBD", x"EDB0", x"EDF9", x"EDA6", x"ED3C", x"ECEA", x"EC10", x"EB3E", x"EB27", x"EAB1", x"E978", x"E8BF", x"E88F", x"E887", x"E981", x"EB50", x"ECA8", x"ED7D", x"EE6D", x"EEEB", x"EECB", x"EEE6", x"EEFE", x"EEF1", x"EF6B", x"F035", x"F0C7", x"F14B", x"F1C8", x"F1D1", x"F1B2", x"F1D5", x"F1C9", x"F1BB", x"F202", x"F1C7", x"F0C0", x"EF7E", x"EE00", x"EC4C", x"EB2B", x"EAA1", x"E9B6", x"E8E6", x"E897", x"E84F", x"E83A", x"E90A", x"E9EE", x"EA5D", x"EAFB", x"EBC9", x"EC20", x"EC8E", x"ED24", x"ECD5", x"EBBB", x"EAB6", x"E9EB", x"E97C", x"EA13", x"EB16", x"EB8D", x"EBAC", x"EBC9", x"EB7C", x"EB0C", x"EAE6", x"EAA3", x"EA5E", x"EA89", x"EB00", x"EB61", x"EBD1", x"EC48", x"EC90", x"ECE0", x"ED3A", x"ED49", x"ED25", x"ED05", x"ECBE", x"EC75", x"EC88", x"ECA0", x"EC99", x"EC96", x"EC84", x"EC37", x"EC06", x"EC19", x"EC2C", x"EC3B", x"EC5A", x"EC69", x"EC77", x"ECB4", x"ECCD", x"ECC1", x"EC9B", x"EC0F", x"EADF", x"E994", x"E87C", x"E78E", x"E76B", x"E83C", x"E920", x"E9A1", x"EA1A", x"EA6C", x"EA05", x"E959", x"E8C2", x"E818", x"E7C1", x"E870", x"E9CB", x"EAE3", x"EB8D", x"EBD0", x"EB9D", x"EB24", x"EAAA", x"EA22", x"E978", x"E8A4", x"E7D4", x"E6FD", x"E5E1", x"E474", x"E32E", x"E23D", x"E177", x"E0ED", x"E102", x"E16E", x"E242", x"E3EF", x"E5F9", x"E76C", x"E88C", x"E9F3", x"EB4F", x"ECB1", x"EE75", x"EF9F", x"EF5F", x"EEB3", x"EE6F", x"EE51", x"EE72", x"EF4F", x"EFCE", x"EF60", x"EEDF", x"EE7C", x"ED89", x"EC4D", x"EB63", x"EA5F", x"E965", x"E908", x"E92A", x"E94D", x"E994", x"EA29", x"EAB5", x"EB29", x"EB8A", x"EBBB", x"EBF4", x"EC57", x"ECF2", x"EDF4", x"EF15", x"EFEF", x"F082", x"F0ED", x"F0AD", x"F014", x"EFA8", x"EF44", x"EE82", x"EE08", x"EDAD", x"ECEB", x"EC97", x"ED65", x"EE59", x"EEDE", x"EF17", x"EE61", x"EC80", x"EB2A", x"EB23", x"EBCA", x"ED00", x"EEDC", x"F020", x"F07E", x"F0A6", x"F04E", x"EF24", x"EDFB", x"ED4B", x"ECC6", x"ECE2", x"EDC5", x"EE7A", x"EECA", x"EEFE", x"EE9B", x"EDD0", x"ED70", x"ED7C", x"ED6D", x"ED7A", x"ED50", x"EC67", x"EB67", x"EB12", x"EAE9", x"EAC8", x"EAFE", x"EAD8", x"EA2C", x"E9E8", x"EA2B", x"EA20", x"EA40", x"EACF", x"EB1C", x"EB4C", x"EC16", x"ECDC", x"ECC9", x"EC60", x"EBB5", x"EA98", x"E9A1", x"E9B9", x"EA4F", x"EB24", x"EC5B", x"ED9D", x"EE6B", x"EEF8", x"EF52", x"EF4B", x"EF63", x"EFF8", x"F0F2", x"F1F8", x"F30A", x"F3AD", x"F3DC", x"F431", x"F4E0", x"F5B6", x"F6A8", x"F775", x"F78B", x"F6DC", x"F605", x"F53C", x"F4B0", x"F4B9", x"F55A", x"F617", x"F72B", x"F8B5", x"FA1B", x"FAC1", x"FAF0", x"FAA1", x"F9E9", x"F9E6", x"FAE0", x"FBE0", x"FC75", x"FD09", x"FD1F", x"FC32", x"FB11", x"FA0B", x"F8A6", x"F7BB", x"F882", x"FA16", x"FB61", x"FC8F", x"FD17", x"FC41", x"FB17", x"FA9E", x"FA49", x"FA34", x"FAE1", x"FB8D", x"FBA9", x"FBF2", x"FC7C", x"FC92", x"FCBA", x"FD20", x"FCCE", x"FC24", x"FC11", x"FBCD", x"FABC", x"F9AF", x"F8B1", x"F774", x"F73C", x"F8A4", x"FA2D", x"FB7D", x"FD0D", x"FE55", x"FED6", x"FFA6", x"0083", x"00BB", x"0104", x"01FB", x"02E6", x"0397", x"0463", x"0449", x"0343", x"0265", x"01D8", x"015D", x"01AC", x"0262", x"0226", x"0144", x"006A", x"FEF2", x"FD5E", x"FCA9", x"FC04", x"FAAF", x"FA04", x"FA58", x"FA8B", x"FB27", x"FC80", x"FD25", x"FD25", x"FE0E", x"FF6B", x"FFF0", x"0024", x"0014", x"FF12", x"FE4B", x"FF37", x"0111", x"02FE", x"0528", x"06D0", x"0761", x"07B3", x"080F", x"07E0", x"076E", x"0719", x"0673", x"05B2", x"0563", x"04F1", x"0403", x"0309", x"0204", x"00BE", x"FFFC", x"002F", x"0105", x"0275", x"0464", x"05C2", x"0623", x"05C6", x"04FE", x"044E", x"047E", x"0551", x"0641", x"075E", x"0860", x"08FC", x"0991", x"0A89", x"0B54", x"0BFA", x"0C86", x"0C49", x"0A9C", x"0833", x"05E0", x"0417", x"03A6", x"04BA", x"0631", x"073F", x"07BD", x"07AD", x"0717", x"069D", x"0674", x"0657", x"0653", x"0666", x"064C", x"05F9", x"05B0", x"0572", x"0515", x"04BA", x"0471", x"0452", x"048D", x"0533", x"061E", x"06E1", x"0751", x"0779", x"078B", x"07D6", x"082F", x"087F", x"08AE", x"089E", x"0887", x"08C5", x"09E4", x"0B79", x"0D30", x"0EDB", x"0FEB", x"0FA0", x"0E39", x"0C57", x"0A4A", x"0890", x"0857", x"0939", x"0A11", x"0ABA", x"0B98", x"0C26", x"0CCF", x"0E45", x"0FBF", x"1035", x"105F", x"10B1", x"10A9", x"10FC", x"1212", x"12F2", x"134C", x"13BD", x"13E7", x"1331", x"129C", x"1241", x"1162", x"106E", x"1007", x"0F70", x"0ECF", x"0EF8", x"0ED5", x"0DAF", x"0CA9", x"0C33", x"0B9F", x"0BD7", x"0D05", x"0DC3", x"0E37", x"0FDA", x"11D3", x"12AB", x"12F5", x"1291", x"10ED", x"0F79", x"0FD1", x"10A1", x"10FB", x"1160", x"1165", x"105F", x"0F63", x"0EEF", x"0E41", x"0D8C", x"0D6A", x"0D42", x"0CBB", x"0C6A", x"0C2D", x"0BCA", x"0C18", x"0CF8", x"0DB3", x"0E7B", x"0F60", x"0FA4", x"0F66", x"0F96", x"0FA4", x"0F77", x"0FC0", x"1033", x"0FC1", x"0F01", x"0E62", x"0D37", x"0BFA", x"0B87", x"0B2C", x"0A73", x"0AB1", x"0BAC", x"0C59", x"0D0A", x"0DBA", x"0CD3", x"0B20", x"0AD6", x"0BCB", x"0D65", x"104E", x"1364", x"147C", x"148C", x"14D3", x"148C", x"13CF", x"13F5", x"1435", x"13BB", x"13CA", x"1493", x"14B6", x"14A5", x"14EA", x"1498", x"13DF", x"13D8", x"13CE", x"1328", x"12CC", x"1288", x"11DB", x"11D6", x"1292", x"12E9", x"130C", x"135B", x"1314", x"1283", x"12E3", x"1340", x"1301", x"1319", x"1360", x"133C", x"140D", x"15E6", x"169E", x"1603", x"151A", x"135E", x"116A", x"1189", x"130A", x"140A", x"14FA", x"163D", x"163D", x"152F", x"1449", x"1290", x"0FCC", x"0DEF", x"0D72", x"0D3E", x"0D60", x"0E26", x"0EA1", x"0F04", x"1027", x"118F", x"124A", x"1271", x"121F", x"1172", x"10FD", x"1161", x"1274", x"140D", x"159E", x"16D2", x"1770", x"178B", x"1755", x"173C", x"173B", x"16EE", x"166F", x"1605", x"15C1", x"15CE", x"166C", x"16EA", x"168B", x"158C", x"147D", x"13EE", x"14B6", x"1743", x"1A92", x"1D74", x"1F72", x"2043", x"1FF3", x"1F1C", x"1E71", x"1E00", x"1DD0", x"1E1C", x"1EC2", x"1F0B", x"1EBC", x"1E4D", x"1E05", x"1DEE", x"1E55", x"1F0F", x"1F3E", x"1E91", x"1D63", x"1BD1", x"198F", x"1760", x"15DC", x"1510", x"1504", x"15AE", x"1676", x"16D3", x"16A9", x"1648", x"15B6", x"1538", x"1504", x"1569", x"164B", x"170B", x"1735", x"16FE", x"1694", x"1671", x"1760", x"197D", x"1B84", x"1D03", x"1DE5", x"1DAD", x"1C2F", x"1A5D", x"1836", x"1581", x"12F5", x"1142", x"0FD8", x"0ECB", x"0E6B", x"0E2A", x"0DBF", x"0DD0", x"0E80", x"0F26", x"0FF4", x"10A9", x"10FA", x"10F7", x"1110", x"114B", x"11D0", x"12AB", x"136C", x"13FE", x"144F", x"13F7", x"1338", x"12B8", x"1224", x"1128", x"1055", x"0FA8", x"0EA8", x"0DAD", x"0CD7", x"0B53", x"092D", x"0786", x"069D", x"06A4", x"0814", x"0A6B", x"0CC9", x"0EED", x"106A", x"10A1", x"1007", x"0F0D", x"0DA2", x"0C31", x"0B2B", x"0A01", x"08D9", x"0893", x"08FD", x"099A", x"0A8E", x"0B68", x"0B52", x"0AB3", x"09F4", x"08D7", x"07EE", x"078C", x"0701", x"064E", x"060C", x"05CD", x"0560", x"05A3", x"05FB", x"056A", x"051A", x"05BE", x"061A", x"062C", x"06E3", x"0746", x"06F4", x"0785", x"08D9", x"093A", x"091B", x"09D9", x"0B0B", x"0CCD", x"0FF1", x"1353", x"1560", x"1643", x"167D", x"15A0", x"13E1", x"11D7", x"0F57", x"0C58", x"0920", x"0618", x"036D", x"018A", x"0072", x"002D", x"006C", x"0073", x"0022", x"FFDF", x"FFAA", x"FF4A", x"FF34", x"FF34", x"FEE0", x"FEA2", x"FF47", x"0053", x"017F", x"0301", x"045D", x"053C", x"0644", x"079A", x"0849", x"083E", x"0803", x"0785", x"06DB", x"06CE", x"06DA", x"0636", x"0571", x"0581", x"0669", x"080D", x"0A90", x"0CE8", x"0E0B", x"0E22", x"0DA2", x"0C53", x"0A77", x"08C7", x"075C", x"0601", x"04DB", x"03F9", x"02EF", x"0195", x"0088", x"0006", x"FFDC", x"0009", x"0070", x"00C7", x"00BC", x"00E3", x"0119", x"00A1", x"FF9B", x"FE9F", x"FDB8", x"FCEA", x"FCFF", x"FD6F", x"FD33", x"FCD1", x"FD1B", x"FD03", x"FC05", x"FB41", x"FAD2", x"FA1D", x"FA2B", x"FB32", x"FB24", x"F97F", x"F836", x"F836", x"F923", x"FBBC", x"FFB9", x"030E", x"04C1", x"058A", x"0509", x"02CA", x"FFAF", x"FCD4", x"FA73", x"F8A2", x"F76C", x"F672", x"F54C", x"F425", x"F351", x"F32A", x"F363", x"F39F", x"F3CF", x"F3DA", x"F3AB", x"F363", x"F349", x"F319", x"F2B3", x"F20C", x"F152", x"F115", x"F1C6", x"F303", x"F452", x"F59C", x"F654", x"F637", x"F641", x"F699", x"F67B", x"F631", x"F68B", x"F69F", x"F5A8", x"F444", x"F24A", x"EF96", x"EE11", x"EF45", x"F239", x"F5CC", x"F956", x"FB5B", x"FB17", x"F9C7", x"F85C", x"F6EF", x"F5F0", x"F5B5", x"F5A0", x"F55E", x"F52D", x"F51A", x"F54A", x"F5CD", x"F65A", x"F69C", x"F65F", x"F563", x"F41E", x"F31D", x"F20C", x"F0CA", x"EFF2", x"EF3B", x"EE66", x"EE49", x"EEEE", x"EF3C", x"EF52", x"EF91", x"EF1E", x"EDF2", x"ED11", x"EC31", x"EB1D", x"EAE8", x"EBBF", x"EC8B", x"ED33", x"ED75", x"EC43", x"EA50", x"E98A", x"EA49", x"EC93", x"F0B7", x"F51F", x"F7E8", x"F8FF", x"F885", x"F5EC", x"F21B", x"EE62", x"EADF", x"E80D", x"E6DD", x"E6EC", x"E771", x"E86E", x"E97D", x"EA51", x"EB39", x"EBFA", x"EC31", x"EC05", x"EB99", x"EAAD", x"EA2A", x"EA52", x"EA6E", x"EA9D", x"EB92", x"EC8F", x"ED5E", x"EEC2", x"F01F", x"F082", x"F0EF", x"F1B6", x"F208", x"F224", x"F2F3", x"F36E", x"F361", x"F385", x"F2EF", x"F0B2", x"EE0C", x"EBFF", x"EAA8", x"EB06", x"ED3C", x"EF69", x"F07C", x"F08E", x"EF3D", x"ECA6", x"EA12", x"E816", x"E67E", x"E5E7", x"E65C", x"E728", x"E83D", x"E9CD", x"EB8E", x"EDA4", x"F04B", x"F2D0", x"F4CD", x"F62D", x"F69D", x"F618", x"F580", x"F4E0", x"F461", x"F498", x"F580", x"F684", x"F7CD", x"F942", x"FA05", x"FA2A", x"FA2C", x"F95C", x"F7BB", x"F656", x"F536", x"F44B", x"F4A5", x"F617", x"F710", x"F769", x"F78A", x"F6FD", x"F67A", x"F78E", x"F9DD", x"FC10", x"FE4D", x"FFF2", x"FFC2", x"FE48", x"FC68", x"F99A", x"F601", x"F314", x"F0E2", x"EF2C", x"EEDD", x"F008", x"F120", x"F219", x"F35C", x"F448", x"F45A", x"F473", x"F48B", x"F3DB", x"F2F7", x"F2CD", x"F2D5", x"F2AF", x"F31C", x"F44F", x"F5AC", x"F729", x"F8E2", x"F9C2", x"F8FC", x"F745", x"F576", x"F366", x"F173", x"F02B", x"EF35", x"EDDA", x"EC58", x"EAE8", x"E90D", x"E779", x"E741", x"E8A4", x"EB0B", x"EE5E", x"F19C", x"F398", x"F465", x"F462", x"F36E", x"F20E", x"F128", x"F08B", x"EFCE", x"EF81", x"EF4A", x"EE7F", x"ED9E", x"ED21", x"EC5D", x"EB82", x"EB26", x"EAC9", x"E9C1", x"E8B7", x"E7A9", x"E640", x"E585", x"E5EA", x"E69A", x"E73B", x"E819", x"E85A", x"E803", x"E83F", x"E8B3", x"E853", x"E7A7", x"E699", x"E4B2", x"E319", x"E33F", x"E421", x"E4EC", x"E606", x"E68C", x"E643", x"E713", x"E9C9", x"ED49", x"F158", x"F5A1", x"F7EB", x"F80B", x"F737", x"F533", x"F20E", x"EF99", x"EDD4", x"EBAD", x"EA2C", x"EA0C", x"E9BF", x"E99A", x"EAC6", x"EC03", x"EC5D", x"ECFF", x"EDBB", x"ED41", x"ECD8", x"ED97", x"EE82", x"EF6E", x"F0F1", x"F23A", x"F2BA", x"F38C", x"F4DC", x"F632", x"F7A8", x"F8E5", x"F933", x"F8BD", x"F7D4", x"F662", x"F539", x"F48F", x"F37C", x"F193", x"EF48", x"EC8D", x"EA6F", x"EAAA", x"ED3D", x"F105", x"F533", x"F8B2", x"FA62", x"FAED", x"FB11", x"FB07", x"FB62", x"FC4B", x"FCA7", x"FC6D", x"FC36", x"FB81", x"FA62", x"FA05", x"F994", x"F870", x"F7F7", x"F8AB", x"F93A", x"F9CF", x"FA90", x"F9E2", x"F7C8", x"F61F", x"F4D7", x"F3A1", x"F39F", x"F489", x"F555", x"F6B8", x"F886", x"F97C", x"F9B5", x"F99B", x"F82A", x"F64E", x"F5B2", x"F537", x"F405", x"F31F", x"F197", x"EEE1", x"EDBB", x"EF99", x"F285", x"F65A", x"FAD2", x"FD18", x"FCA3", x"FBD0", x"FA9D", x"F8A7", x"F7B9", x"F77E", x"F5F9", x"F459", x"F3D0", x"F34A", x"F3BA", x"F63F", x"F885", x"F987", x"FAF5", x"FC39", x"FC4F", x"FD12", x"FE3E", x"FDA3", x"FC4A", x"FBEA", x"FB19", x"FA23", x"FA9B", x"FB3D", x"FB26", x"FC17", x"FDC3", x"FEB9", x"FF9D", x"0059", x"FF48", x"FD8D", x"FC6D", x"FADE", x"F8DE", x"F761", x"F516", x"F217", x"F0F6", x"F233", x"F4E6", x"F9A4", x"FF23", x"0282", x"03DB", x"0424", x"02A9", x"0051", x"FEDB", x"FD64", x"FB89", x"FA97", x"FA19", x"F934", x"F910", x"F97C", x"F929", x"F8EE", x"F95E", x"F95C", x"F973", x"FA56", x"FA7C", x"F9B6", x"F924", x"F824", x"F6E9", x"F79E", x"F9A4", x"FB41", x"FD64", x"FF7F", x"FF79", x"FF27", x"002B", x"000B", x"FED6", x"FF28", x"FFF9", x"0032", x"0243", x"04E7", x"0486", x"02B5", x"027A", x"02BA", x"0466", x"08F5", x"0D60", x"0EF1", x"0F4E", x"0E74", x"0B62", x"0830", x"05BA", x"0279", x"FF48", x"FD21", x"FAB8", x"F8AB", x"F8EA", x"FA25", x"FB52", x"FD95", x"FF98", x"000E", x"00DA", x"0236", x"0227", x"0192", x"01D7", x"018F", x"014C", x"027F", x"03A5", x"03AF", x"0428", x"0490", x"03D3", x"030D", x"020C", x"FF45", x"FC09", x"F9C5", x"F7D0", x"F73B", x"F90A", x"FAA0", x"FA74", x"F9C3", x"F87F", x"F70F", x"F88F", x"FD14", x"0196", x"0559", x"0872", x"094F", x"08B8", x"08DB", x"0903", x"085A", x"07E8", x"07A4", x"06E3", x"0690", x"06D2", x"0714", x"07B9", x"08BB", x"0941", x"09FF", x"0B0F", x"0B78", x"0BFB", x"0CFA", x"0CAC", x"0B41", x"0A96", x"09DF", x"08AC", x"08E1", x"0985", x"086E", x"073E", x"06CD", x"0540", x"033F", x"0285", x"0156", x"0010", x"01A4", x"0501", x"07A0", x"0A27", x"0B76", x"0967", x"06FA", x"0769", x"0901", x"0B32", x"0EAE", x"1064", x"0ED0", x"0D28", x"0C4F", x"0AA0", x"0958", x"0920", x"07A9", x"0598", x"04EF", x"04F7", x"051F", x"06C1", x"08DD", x"0A17", x"0B38", x"0C1A", x"0BEC", x"0BAE", x"0BDD", x"0B9C", x"0B5A", x"0BB6", x"0BBF", x"0B47", x"0ACA", x"0998", x"07DF", x"069D", x"0585", x"0489", x"0439", x"03BF", x"02C9", x"02B0", x"0307", x"02C8", x"033F", x"0405", x"0266", x"FF56", x"FD23", x"FB53", x"FAE1", x"FE86", x"03BF", x"06F4", x"0915", x"0AD7", x"0AB2", x"0A70", x"0BE6", x"0C80", x"0B5B", x"0A52", x"0904", x"067F", x"04F4", x"0494", x"0403", x"042E", x"058D", x"066D", x"06E2", x"07AC", x"07B4", x"0735", x"07A6", x"0897", x"0935", x"0A18", x"0A3A", x"08E4", x"0796", x"06CB", x"05F6", x"05E9", x"068F", x"062D", x"05A8", x"05D1", x"056C", x"0503", x"0688", x"0810", x"079E", x"0689", x"0479", x"00B8", x"FEBC", x"0099", x"035A", x"05C4", x"08B3", x"0A39", x"09C2", x"09E6", x"0A97", x"09BF", x"0897", x"07F1", x"06BF", x"0573", x"0580", x"0603", x"06DB", x"08B8", x"0A82", x"0B86", x"0C7B", x"0D34", x"0D90", x"0E82", x"0F9B", x"0FA4", x"0F68", x"0F0C", x"0D8D", x"0BCF", x"0AA8", x"0907", x"0747", x"06B2", x"0657", x"05BD", x"0616", x"0672", x"0612", x"0694", x"0838", x"095C", x"0AAB", x"0BEF", x"0B2E", x"09B0", x"0A65", x"0C6B", x"0EF5", x"130D", x"167E", x"16FC", x"1723", x"1847", x"183B", x"17C3", x"17FD", x"16F1", x"14BE", x"1496", x"15C0", x"164E", x"1732", x"1820", x"1755", x"164D", x"166D", x"163F", x"15A2", x"157E", x"148B", x"1280", x"10C9", x"0F03", x"0CD0", x"0BB3", x"0B34", x"0A50", x"0A3D", x"0B2A", x"0BF1", x"0DB3", x"10DC", x"1328", x"14D4", x"1793", x"19B3", x"1A75", x"1B7D", x"1B26", x"1794", x"140F", x"1301", x"12A0", x"13E6", x"177F", x"194B", x"17EF", x"16DE", x"16A6", x"15DA", x"1681", x"18D8", x"19B6", x"1959", x"1998", x"191F", x"1749", x"1610", x"15D2", x"15CC", x"164C", x"16D3", x"163E", x"1507", x"13B6", x"126B", x"119C", x"10A6", x"0ED3", x"0D4E", x"0CA5", x"0B64", x"0A16", x"09C1", x"0925", x"088A", x"0995", x"0AEB", x"0ACE", x"0AF2", x"0BCB", x"0C03", x"0CA4", x"0DE9", x"0D09", x"0A22", x"0752", x"04A0", x"030C", x"0533", x"091C", x"0B78", x"0C9E", x"0C8B", x"0A17", x"088B", x"0A0B", x"0B73", x"0B47", x"0B12", x"092A", x"04C5", x"01A5", x"0028", x"FE0E", x"FCB3", x"FD66", x"FD8D", x"FD3F", x"FE79", x"FF9C", x"FFAE", x"006B", x"0110", x"0028", x"FF78", x"FF6E", x"FE6E", x"FDB4", x"FE70", x"FEE1", x"FF1D", x"0096", x"0178", x"00D1", x"0171", x"03CD", x"05F5", x"081D", x"09DA", x"08A4", x"0517", x"02B9", x"0277", x"03AD", x"0680", x"09FF", x"0C58", x"0D55", x"0DCA", x"0DDB", x"0D78", x"0CEA", x"0D23", x"0E0B", x"0E6B", x"0D99", x"0C3E", x"0A4E", x"0831", x"07AA", x"0857", x"0800", x"0708", x"069E", x"0604", x"05C6", x"0724", x"080D", x"06D5", x"05BC", x"051E", x"0369", x"0228", x"01E9", x"FFC1", x"FC8E", x"FBE4", x"FC9B", x"FD01", x"FF40", x"027D", x"03A9", x"0502", x"085A", x"0A18", x"0918", x"0847", x"0790", x"06DD", x"09A5", x"0F7A", x"13FE", x"1626", x"1702", x"1588", x"12C1", x"1175", x"1120", x"1058", x"0FE6", x"0F6F", x"0DEE", x"0C56", x"0B75", x"0A7C", x"098D", x"091C", x"087C", x"07EF", x"08AE", x"0A5B", x"0C42", x"0E34", x"0F36", x"0E53", x"0CA6", x"0B5C", x"0AB2", x"0B3F", x"0D1F", x"0EC6", x"0F45", x"0F04", x"0E59", x"0D70", x"0D5F", x"0F1B", x"11B1", x"13CE", x"14BB", x"13ED", x"10C6", x"0CC0", x"0A47", x"097A", x"093B", x"0A03", x"0C37", x"0E0A", x"0F29", x"1073", x"1036", x"0D26", x"0A0B", x"08E0", x"07AC", x"067D", x"068C", x"0614", x"0435", x"038D", x"040F", x"030C", x"0154", x"0072", x"FF31", x"FDEF", x"FE9B", x"000D", x"0095", x"013B", x"01E8", x"0197", x"0163", x"0211", x"01FF", x"0143", x"0115", x"0111", x"0169", x"0398", x"069F", x"090A", x"0B7D", x"0E4D", x"100E", x"1073", x"0FDB", x"0E16", x"0BE0", x"0B00", x"0BE3", x"0DB0", x"0FAD", x"111F", x"121C", x"129A", x"121D", x"10E1", x"101B", x"0F9C", x"0EFA", x"0EF0", x"0EBD", x"0CCA", x"0A4A", x"0915", x"083F", x"06FF", x"05E8", x"0471", x"01C6", x"FF9B", x"FF42", x"FFFA", x"0149", x"0328", x"0491", x"04CA", x"03EF", x"0269", x"00D5", x"FFD2", x"FF14", x"FE8C", x"FE48", x"FD8B", x"FC98", x"FC6C", x"FD02", x"FD5C", x"FDC1", x"FDAC", x"FC11", x"F98F", x"F75B", x"F5BA", x"F5A3", x"F807", x"FBD7", x"FFFF", x"045D", x"0712", x"0707", x"059F", x"0404", x"0236", x"01D8", x"0322", x"0363", x"01B4", x"FFD0", x"FDBE", x"FBD8", x"FB79", x"FB9F", x"FA36", x"F825", x"F65F", x"F4C7", x"F498", x"F615", x"F6D5", x"F640", x"F54C", x"F30D", x"F054", x"EFD9", x"F07E", x"EF39", x"ED4D", x"EBCA", x"E98D", x"E86D", x"EAC1", x"EDCF", x"EF5B", x"F114", x"F2E2", x"F2BE", x"F14D", x"EFFF", x"EEE6", x"EEDF", x"F0DD", x"F3EC", x"F692", x"F7E7", x"F7FE", x"F87E", x"F93D", x"F884", x"F784", x"F828", x"F83E", x"F6CD", x"F5CB", x"F403", x"F01A", x"EED0", x"F22A", x"F50E", x"F5E1", x"F6A5", x"F547", x"F17F", x"F091", x"F24D", x"F1DC", x"F04D", x"EF7F", x"ECCC", x"E931", x"E88D", x"E901", x"E7EF", x"E82F", x"EA0E", x"EAFE", x"EBFD", x"EE7C", x"EFC6", x"EFB9", x"F165", x"F443", x"F5B1", x"F597", x"F477", x"F22D", x"F061", x"F13F", x"F44D", x"F6EE", x"F802", x"F8C1", x"F9B3", x"F9A8", x"F8F6", x"F8FF", x"F8A2", x"F72A", x"F6D4", x"F721", x"F508", x"F22B", x"F1FF", x"F2D8", x"F333", x"F494", x"F4FD", x"F231", x"EF94", x"EFA1", x"EFD5", x"EFFD", x"F0FB", x"F023", x"ECEB", x"EABA", x"E96D", x"E7AE", x"E759", x"E863", x"E85C", x"E909", x"EC50", x"EF72", x"F18A", x"F407", x"F564", x"F47C", x"F41B", x"F47E", x"F355", x"F175", x"F0B7", x"F07D", x"F0E6", x"F27F", x"F3A8", x"F347", x"F1EA", x"EFDE", x"EE21", x"EDF4", x"EE7B", x"EF5E", x"F0EB", x"F111", x"EE0A", x"EA8E", x"E867", x"E68B", x"E5FB", x"E754", x"E6EA", x"E3B8", x"E1AD", x"E11B", x"DFEA", x"DF1A", x"DECF", x"DC5C", x"D93A", x"D8C1", x"D9E9", x"DAF2", x"DCFA", x"DEC2", x"DE24", x"DD01", x"DD29", x"DD65", x"DE1C", x"E09E", x"E300", x"E383", x"E39A", x"E362", x"E191", x"DFD8", x"E083", x"E2F6", x"E67D", x"EB6E", x"EFEF", x"F1A5", x"F192", x"F140", x"F0E3", x"F09F", x"F141", x"F1F4", x"F1EB", x"F10E", x"EF46", x"ED06", x"EB77", x"EAE9", x"EAD6", x"EB2A", x"EAC7", x"E8C9", x"E723", x"E733", x"E746", x"E6B3", x"E6FB", x"E6EC", x"E532", x"E3D2", x"E300", x"E075", x"DDE6", x"DE45", x"DF7C", x"DFB2", x"E046", x"E0C5", x"E023", x"E10C", x"E448", x"E6DC", x"E838", x"E92A", x"E885", x"E701", x"E72D", x"E891", x"EAD0", x"EF02", x"F2D6", x"F39F", x"F33E", x"F29E", x"F09F", x"EFB4", x"F109", x"F11C", x"F021", x"F1A2", x"F396", x"F3AE", x"F45E", x"F4DC", x"F269", x"F086", x"F1CC", x"F248", x"F13A", x"F122", x"F050", x"EE51", x"EEC4", x"F0CF", x"F080", x"EE9F", x"EBE8", x"E746", x"E333", x"E2A4", x"E3C3", x"E597", x"E861", x"E97C", x"E812", x"E6E0", x"E64D", x"E5AC", x"E66E", x"E75A", x"E587", x"E247", x"DFC2", x"DDBC", x"DD7A", x"E04D", x"E347", x"E491", x"E4E9", x"E351", x"DF90", x"DC4D", x"DA11", x"D867", x"D913", x"DBBD", x"DDCA", x"DF84", x"E0E0", x"DFC2", x"DD4F", x"DC24", x"DB0F", x"DA26", x"DB4D", x"DCE2", x"DCC0", x"DCEA", x"DD36", x"DC16", x"DBC5", x"DD58", x"DE46", x"DEE9", x"E046", x"E08C", x"E02A", x"E21B", x"E481", x"E5CA", x"E7A7", x"E95D", x"E997", x"EB7A", x"EEEA", x"F035", x"F009", x"EFB5", x"ED5A", x"EB1C", x"ECD8", x"EFC1", x"F1A6", x"F4A2", x"F68B", x"F4AC", x"F326", x"F360", x"F1D9", x"F034", x"F0E4", x"F04D", x"EE6B", x"EEDA", x"EF4E", x"ED4C", x"EBDB", x"EB2E", x"E8E4", x"E74E", x"E76D", x"E654", x"E4EF", x"E4D6", x"E3E3", x"E2A6", x"E3BB", x"E53E", x"E681", x"E99B", x"EBE0", x"EB01", x"EABF", x"EBB0", x"EAE6", x"EAE0", x"ED05", x"ED80", x"ED76", x"F08B", x"F2F6", x"F1E0", x"F0C3", x"EF6C", x"EC2B", x"EB45", x"EE05", x"EFC0", x"F093", x"F2C5", x"F3CE", x"F364", x"F463", x"F53B", x"F3E1", x"F2BD", x"F275", x"F1C4", x"F23E", x"F43E", x"F5AB", x"F69A", x"F76B", x"F6F8", x"F682", x"F774", x"F878", x"F9F6", x"FCB3", x"FD72", x"FB61", x"F9A1", x"F7EF", x"F580", x"F5AA", x"F7BE", x"F73F", x"F619", x"F7C5", x"F9A9", x"FB33", x"FEBB", x"012E", x"FFEF", x"FF43", x"00C3", x"0156", x"0149", x"01EE", x"012A", x"FF74", x"FFCE", x"016C", x"02A5", x"0411", x"0578", x"0639", x"0741", x"089D", x"0A00", x"0C20", x"0E03", x"0E42", x"0DEF", x"0D89", x"0CAB", x"0D67", x"1055", x"11C2", x"10BE", x"0F57", x"0D81", x"0C34", x"0ED5", x"13CE", x"16CF", x"1817", x"183F", x"1609", x"13FC", x"1509", x"168E", x"16F7", x"1801", x"18BD", x"17F4", x"183B", x"1994", x"188A", x"15D1", x"13C5", x"11DA", x"10AC", x"1217", x"144D", x"14DB", x"1477", x"13DB", x"12B4", x"122C", x"12E8", x"146C", x"1680", x"1807", x"17C6", x"16C6", x"15ED", x"14CF", x"1497", x"15DF", x"15F9", x"1480", x"1472", x"1590", x"15C5", x"1658", x"17B9", x"1770", x"166D", x"172C", x"17D1", x"1667", x"14C0", x"1351", x"10F4", x"0EFA", x"0E54", x"0D89", x"0C68", x"0C01", x"0BC3", x"0B9C", x"0C9B", x"0E83", x"1040", x"1235", x"13D2", x"143E", x"148B", x"156D", x"161F", x"1668", x"1735", x"17DE", x"1808", x"187B", x"192B", x"19B7", x"1ADF", x"1CA7", x"1DF8", x"1E46", x"1D83", x"1B84", x"193F", x"17C8", x"16B0", x"1576", x"14A5", x"13BD", x"1228", x"10BD", x"1011", x"0F81", x"0F44", x"0FBC", x"0FEB", x"0F0B", x"0DA7", x"0C00", x"0A89", x"0A24", x"0AFB", x"0CBB", x"0F30", x"1189", x"12E2", x"145C", x"165B", x"17C3", x"18B6", x"1A13", x"1A8A", x"1A1D", x"1AB2", x"1B7B", x"199B", x"163E", x"137D", x"1136", x"1038", x"1213", x"1426", x"137C", x"116C", x"0FB1", x"0DBA", x"0C66", x"0CD3", x"0D4F", x"0CC6", x"0C36", x"0BBA", x"0A94", x"09A7", x"09D0", x"0AA8", x"0B75", x"0BB8", x"0AF4", x"09A0", x"08DE", x"0984", x"0BD3", x"0E24", x"0ECB", x"0DE8", x"0C65", x"0A8C", x"0953", x"09BD", x"0AB8", x"0B67", x"0C95", x"0E07", x"0E83", x"0ED6", x"1083", x"1374", x"175C", x"1BDB", x"1F60", x"206A", x"1F3A", x"1D07", x"1B03", x"19DB", x"1A0A", x"1C2A", x"1FCC", x"22C8", x"23FC", x"2388", x"213D", x"1E1D", x"1D27", x"1E53", x"1F18", x"1F2F", x"1F16", x"1D8A", x"1BD8", x"1C74", x"1DBC", x"1D94", x"1D28", x"1C35", x"1973", x"1718", x"16E5", x"16D2", x"16C2", x"1838", x"1950", x"1899", x"17AA", x"165A", x"13AE", x"11AC", x"10F6", x"0FF4", x"0E98", x"0D5F", x"0BB0", x"0A8C", x"0B1F", x"0BB8", x"0BAA", x"0B35", x"0871", x"033A", x"FE9C", x"FB4C", x"F93D", x"FB0A", x"FFD5", x"02E7", x"0397", x"0362", x"0135", x"FEAA", x"FF34", x"0122", x"0208", x"037A", x"0545", x"05FA", x"07B7", x"0AD0", x"0CBA", x"0DC4", x"0EA7", x"0D69", x"0BB8", x"0CE5", x"0EF9", x"106D", x"12D7", x"13AB", x"1111", x"0FA5", x"10B6", x"1002", x"0EE8", x"0FCB", x"0F76", x"0E78", x"1139", x"1479", x"1434", x"14A8", x"174A", x"18CD", x"1ADB", x"1EA9", x"1F42", x"1C92", x"1BDF", x"1D11", x"1ED5", x"2397", x"292F", x"2B29", x"2A91", x"28FF", x"250F", x"2189", x"216E", x"21B0", x"2078", x"1F49", x"1C89", x"1788", x"146B", x"13EF", x"12D2", x"1217", x"134E", x"138F", x"124F", x"11BE", x"10C0", x"0E34", x"0CB0", x"0CCF", x"0C3C", x"0AEA", x"09C1", x"0878", x"07E3", x"08F9", x"0A35", x"0A8E", x"0A24", x"0849", x"05A4", x"04BB", x"05CD", x"07AC", x"0AAD", x"0D5F", x"0C40", x"080E", x"04C0", x"0313", x"030E", x"0620", x"0A38", x"0B15", x"09C5", x"0940", x"0814", x"05F7", x"0515", x"045A", x"01A0", x"0023", x"01AE", x"034D", x"04BB", x"07D7", x"09C1", x"08A7", x"07AC", x"067D", x"023A", x"FE18", x"FDB3", x"FEB6", x"008F", x"04AE", x"0722", x"04C4", x"01B5", x"005A", x"FEB1", x"FDEC", x"FF35", x"FF68", x"FE59", x"FEF6", x"0033", x"0078", x"012D", x"01DF", x"00F3", x"FFF9", x"FF3C", x"FD56", x"FC16", x"FCCE", x"FD59", x"FDFA", x"0033", x"0200", x"02CF", x"04E8", x"065E", x"047C", x"0241", x"019B", x"0077", x"0020", x"01CC", x"020C", x"004C", x"00D0", x"035B", x"04B2", x"056F", x"0533", x"0199", x"FCDF", x"FB8B", x"FD11", x"FF67", x"02DB", x"06E9", x"0984", x"0AD9", x"0C8A", x"0E43", x"0EE8", x"0F09", x"0FBB", x"0F6E", x"0C59", x"0885", x"05FB", x"041D", x"039D", x"05BE", x"071B", x"0512", x"02A1", x"01A9", x"00AD", x"0153", x"0447", x"057E", x"04D7", x"061F", x"088C", x"0A50", x"0D79", x"0FCE", x"0D60", x"09B0", x"0850", x"06EA", x"0668", x"0923", x"0B24", x"0AB7", x"0C38", x"0F0B", x"0F1A", x"0DD2", x"0BD7", x"0680", x"0090", x"FE64", x"FE13", x"FE6F", x"0094", x"01D2", x"008D", x"FFB4", x"FF2C", x"FDA3", x"FD29", x"FD4C", x"FB46", x"F9A6", x"FAE0", x"FC9D", x"FF3C", x"03A0", x"04F2", x"019E", x"FE6E", x"FC55", x"FACE", x"FD7C", x"0325", x"05E1", x"06A8", x"081F", x"07A7", x"0654", x"07A4", x"0869", x"05E4", x"0437", x"0345", x"0005", x"FD31", x"FC85", x"FAB4", x"F8F2", x"FA42", x"FB79", x"FA81", x"F99C", x"F82B", x"F546", x"F44A", x"F603", x"F78E", x"F926", x"FB10", x"FB63", x"FAFC", x"FBFD", x"FD14", x"FD76", x"FE00", x"FDD7", x"FCC3", x"FC9C", x"FD72", x"FE5D", x"FFE7", x"0137", x"00F1", x"0052", x"FF97", x"FDE9", x"FD86", x"FF90", x"012C", x"01A9", x"020F", x"004E", x"FC64", x"FA2D", x"F9AD", x"F831", x"F74F", x"F81A", x"F82A", x"F782", x"F7AF", x"F70F", x"F54B", x"F525", x"F72F", x"F9F3", x"FC8E", x"FDCD", x"FD0B", x"FB79", x"FA05", x"F936", x"FA41", x"FC8F", x"FEFF", x"025F", x"056A", x"0539", x"031D", x"01DE", x"00B5", x"0095", x"0362", x"05E4", x"0597", x"05EE", x"07A4", x"07F3", x"084F", x"09AF", x"089B", x"066C", x"077B", x"09FD", x"0B60", x"0D5E", x"0E9B", x"0C7C", x"0A26", x"09C0", x"08EB", x"083F", x"0969", x"0A03", x"09AD", x"0AA6", x"0B57", x"0A53", x"09AD", x"0968", x"082C", x"0851", x"09B6", x"09A8", x"089A", x"07B2", x"04E8", x"019F", x"00C6", x"00DA", x"0140", x"03B9", x"0508", x"01FA", x"FDF7", x"FA90", x"F665", x"F471", x"F5C7", x"F4D6", x"F182", x"F0D5", x"F14B", x"F04B", x"F091", x"F08A", x"EC0A", x"E7A7", x"E83C", x"EA1C", x"EBD0", x"EF2F", x"F0CB", x"EE97", x"ED51", x"EE54", x"EE63", x"EF06", x"F186", x"F268", x"F1B5", x"F24D", x"F278", x"F096", x"EFA8", x"F076", x"F11C", x"F2B3", x"F5AA", x"F6AC", x"F4BA", x"F2AF", x"F173", x"F069", x"F029", x"F0AF", x"F0AA", x"EFD8", x"EFA1", x"F048", x"F049", x"EF3F", x"EEAC", x"EF52", x"F022", x"F136", x"F304", x"F422", x"F450", x"F58A", x"F728", x"F6F7", x"F5CD", x"F540", x"F4D1", x"F5E3", x"FA01", x"FE9A", x"00FF", x"01C7", x"0067", x"FC2B", x"F83B", x"F6A9", x"F59A", x"F4CB", x"F542", x"F4CA", x"F221", x"EF47", x"EC60", x"E890", x"E5D6", x"E5A5", x"E65C", x"E72E", x"E7B6", x"E63C", x"E2F0", x"DF90", x"DCA4", x"DB0B", x"DBDE", x"DD8D", x"DE7D", x"DF7E", x"E008", x"DF27", x"DEF2", x"E010", x"E005", x"DEE8", x"DEE8", x"DF45", x"DFA6", x"E1AE", x"E3F0", x"E402", x"E369", x"E3A3", x"E433", x"E5FA", x"E96D", x"EBF3", x"ECA4", x"EC8B", x"EAFF", x"E877", x"E791", x"E7D7", x"E77C", x"E778", x"E7C0", x"E69E", x"E5A0", x"E67F", x"E745", x"E763", x"E87D", x"E9D7", x"EA4C", x"EB59", x"EC4A", x"EAE7", x"E828", x"E555", x"E23C", x"E077", x"E1AC", x"E495", x"E826", x"EC2A", x"EE74", x"EDB6", x"EBD1", x"E969", x"E6E5", x"E675", x"E84D", x"EA5E", x"ECB5", x"EF27", x"EF5D", x"ED6F", x"EB56", x"E8DE", x"E71B", x"E8EE", x"ED52", x"F172", x"F538", x"F781", x"F621", x"F34B", x"F19A", x"F015", x"EF44", x"F09C", x"F243", x"F293", x"F36F", x"F453", x"F3D9", x"F3D4", x"F51A", x"F5DB", x"F6E5", x"F8CB", x"F942", x"F7B4", x"F597", x"F1FA", x"ED4E", x"EAAF", x"EA61", x"EB78", x"EEF7", x"F330", x"F465", x"F3A4", x"F2B2", x"F0C2", x"EF82", x"F15A", x"F345", x"F362", x"F447", x"F506", x"F325", x"F128", x"F07D", x"EF08", x"EE91", x"F1EF", x"F5B6", x"F769", x"F8D0", x"F904", x"F67E", x"F48C", x"F430", x"F2EC", x"F15E", x"F160", x"F11B", x"F088", x"F1CD", x"F366", x"F348", x"F36D", x"F48E", x"F59A", x"F78E", x"FA8F", x"FBA4", x"F9C3", x"F6A1", x"F30A", x"EF70", x"ED3A", x"EC9D", x"ED19", x"EED3", x"F122", x"F332", x"F451", x"F3D6", x"F236", x"F141", x"F0F8", x"F075", x"F0B4", x"F218", x"F2E4", x"F2C4", x"F22B", x"EFB9", x"EC09", x"EA81", x"EC2C", x"EFC0", x"F4DC", x"F9DD", x"FC08", x"FBD6", x"FB1A", x"F978", x"F7C4", x"F736", x"F66D", x"F487", x"F39C", x"F435", x"F531", x"F73A", x"FA26", x"FB7C", x"FB12", x"FABD", x"F9F2", x"F84E", x"F6DD", x"F5A4", x"F3AF", x"F198", x"EFB2", x"EE65", x"EF18", x"F18C", x"F3EB", x"F597", x"F5B0", x"F343", x"F0DA", x"F104", x"F191", x"F131", x"F1DC", x"F2B3", x"F189", x"F08C", x"EFF9", x"EC97", x"E850", x"E7E9", x"EA6A", x"EDBF", x"F2B6", x"F6D0", x"F658", x"F40C", x"F2B8", x"F0E9", x"EF09", x"EED4", x"EDD6", x"EB3E", x"E9F3", x"EA0C", x"EA12", x"EBA8", x"EE8C", x"F00D", x"F11D", x"F2F6", x"F3B1", x"F342", x"F3CA", x"F37E", x"F1B4", x"F0D3", x"F0A8", x"F014", x"F167", x"F51A", x"F843", x"FB2C", x"FE9D", x"FFA8", x"FE30", x"FCE7", x"FAF5", x"F864", x"F8B5", x"FB70", x"FCEE", x"FD9E", x"FDA8", x"FAD0", x"F7E7", x"F8CA", x"FB60", x"FDB3", x"011A", x"0381", x"02E9", x"02DA", x"0491", x"04C4", x"03D9", x"0336", x"00F4", x"FD94", x"FCB6", x"FD3B", x"FCCB", x"FC73", x"FC50", x"FB64", x"FB81", x"FD68", x"FEF0", x"FF38", x"FE6E", x"FBAD", x"F7DF", x"F522", x"F317", x"F1F2", x"F2DA", x"F497", x"F59A", x"F6E7", x"F7D1", x"F6A1", x"F482", x"F222", x"EE7E", x"EB2A", x"EA4D", x"EACD", x"EBD9", x"EDAE", x"EDE5", x"EB97", x"E979", x"E8AA", x"E8B9", x"EB06", x"EEE0", x"F10E", x"F17D", x"F1B4", x"F0BD", x"EEE0", x"EE2D", x"EDFF", x"ED60", x"EDB6", x"EED8", x"EFBE", x"F167", x"F3AD", x"F552", x"F719", x"F923", x"FA1D", x"FB57", x"FDE6", x"FF33", x"FEA6", x"FE5C", x"FD4B", x"FB39", x"FBAF", x"FE64", x"FFA8", x"0095", x"0264", x"02C0", x"02AF", x"04DA", x"068D", x"05BF", x"0520", x"049F", x"0347", x"0459", x"07D0", x"08A9", x"070E", x"05AD", x"0399", x"021F", x"055D", x"0A4B", x"0C4A", x"0DA6", x"1013", x"10DC", x"110A", x"12BB", x"1330", x"113B", x"103E", x"1074", x"0FBB", x"0EDD", x"0F37", x"1004", x"115B", x"12D8", x"1376", x"1330", x"124C", x"1055", x"0E43", x"0C17", x"0834", x"0416", x"0321", x"03B3", x"0406", x"064C", x"09E0", x"0B6C", x"0C2E", x"0DA9", x"0BE3", x"06E9", x"0444", x"0489", x"04E5", x"0698", x"08B3", x"06C7", x"0284", x"017F", x"02E8", x"0473", x"0748", x"09D4", x"08EE", x"073F", x"0819", x"0945", x"0961", x"0A07", x"0A3B", x"0844", x"05FF", x"04A3", x"02CE", x"0111", x"01C7", x"0484", x"070E", x"0863", x"0844", x"0674", x"038F", x"0182", x"0114", x"00B9", x"FF6C", x"FEC7", x"FF2D", x"FEBC", x"FDE6", x"FE7E", x"FF30", x"FF79", x"01D6", x"051E", x"04DD", x"0260", x"013A", x"006A", x"FF6E", x"00A0", x"0196", x"FEFD", x"FC98", x"FE37", x"019D", x"055B", x"0A25", x"0D3B", x"0CFB", x"0C4B", x"0C9F", x"0C1C", x"0B4B", x"0B3E", x"0B7A", x"0B81", x"0B61", x"0ACB", x"0A25", x"0A24", x"0AAE", x"0C22", x"0E44", x"0F86", x"10AC", x"1339", x"1556", x"1552", x"1481", x"1246", x"0DFD", x"0B2F", x"0B92", x"0C61", x"0DCD", x"110D", x"133F", x"13CD", x"15E1", x"17C7", x"16A6", x"1579", x"1597", x"1483", x"1437", x"1691", x"171D", x"14E6", x"1488", x"1610", x"17B6", x"1BA7", x"20B9", x"22BA", x"2331", x"24DB", x"257E", x"243E", x"229F", x"1F0B", x"19A5", x"1609", x"145F", x"1361", x"143A", x"161E", x"1672", x"16D2", x"186D", x"1962", x"1A7A", x"1D54", x"1EB0", x"1D4B", x"1C05", x"1A90", x"17DE", x"166E", x"165B", x"14E1", x"13D6", x"157E", x"1819", x"1B09", x"1EC4", x"204D", x"1E3E", x"1B4E", x"1880", x"159B", x"14B1", x"151B", x"142D", x"12A7", x"123E", x"1260", x"1444", x"18CF", x"1D12", x"1F25", x"2009", x"1F0A", x"1C48", x"1A87", x"19D3", x"1850", x"16F0", x"15D3", x"133F", x"10E1", x"10E9", x"1160", x"11B6", x"133B", x"1465", x"1450", x"1593", x"17B9", x"17ED", x"169E", x"148D", x"1061", x"0BF1", x"09FF", x"0971", x"0983", x"0B76", x"0DFF", x"0FC4", x"11F1", x"13FD", x"1442", x"13A6", x"12D8", x"10C8", x"0EBA", x"0DD1", x"0C70", x"0AA8", x"0A28", x"0A14", x"0A46", x"0CBC", x"1036", x"12AB", x"1507", x"16F4", x"1653", x"146D", x"1307", x"10C4", x"0E96", x"0E5A", x"0E0E", x"0C7E", x"0C1D", x"0C63", x"0BE0", x"0CAD", x"0EC3", x"0F2F", x"0F4B", x"10EF", x"114C", x"0FD2", x"0F7D", x"0F49", x"0E4F", x"0FD5", x"1359", x"14DC", x"1538", x"164B", x"1643", x"1615", x"1879", x"1B1A", x"1BDC", x"1CC3", x"1D98", x"1CA2", x"1BEF", x"1BC9", x"1917", x"14BB", x"1194", x"0F91", x"0FD9", x"14C8", x"1B14", x"1EB7", x"2086", x"2134", x"2007", x"1F50", x"203F", x"1FDE", x"1D70", x"1B0C", x"1861", x"15AD", x"150C", x"1611", x"1707", x"1862", x"1971", x"187B", x"16DA", x"15D5", x"1404", x"116C", x"0F4B", x"0C72", x"090C", x"0810", x"0948", x"0A43", x"0B6C", x"0D48", x"0DF6", x"0D9D", x"0DA2", x"0D04", x"0B06", x"0923", x"0803", x"06BD", x"0545", x"03B0", x"01AD", x"FF5D", x"FD43", x"FBB2", x"FB7C", x"FCCE", x"FEE1", x"0166", x"038F", x"045B", x"0424", x"0444", x"049D", x"047D", x"0433", x"0378", x"01D4", x"FFFF", x"FEC6", x"FE25", x"FE5A", x"FF8B", x"0133", x"02C0", x"03F9", x"0510", x"0684", x"0875", x"0A00", x"0AB5", x"0A50", x"0891", x"06D4", x"06F8", x"0856", x"09EF", x"0BDA", x"0CA1", x"0B08", x"095B", x"0970", x"0967", x"094B", x"0A7E", x"0AE5", x"0930", x"082A", x"0800", x"05D9", x"039A", x"042F", x"05EB", x"075A", x"0A28", x"0C7C", x"0BBF", x"0A55", x"0AB3", x"0B0C", x"0A72", x"0A64", x"0A94", x"0A42", x"0A7D", x"0B9F", x"0C15", x"0B3A", x"09FF", x"0924", x"0827", x"0649", x"046B", x"0395", x"0357", x"035A", x"03FB", x"0365", x"FFCD", x"FBA1", x"F94A", x"F779", x"F600", x"F667", x"F703", x"F64E", x"F6F5", x"F970", x"FA60", x"FA2E", x"FB4A", x"FBF5", x"FAF9", x"FAD0", x"FA89", x"F79E", x"F4EF", x"F5AF", x"F7BD", x"F9F8", x"FD63", x"FF96", x"FE79", x"FD52", x"FDC6", x"FD7E", x"FC8E", x"FC51", x"FB03", x"F85C", x"F749", x"F7BA", x"F78F", x"F77D", x"F832", x"F815", x"F73C", x"F73A", x"F70E", x"F5CF", x"F4A8", x"F3E6", x"F2B6", x"F1A4", x"F11A", x"F0E2", x"F127", x"F22B", x"F31F", x"F3DC", x"F420", x"F36C", x"F26B", x"F278", x"F2F0", x"F432", x"F7AC", x"FBC2", x"FDA1", x"FD4C", x"FB06", x"F675", x"F2C2", x"F3BD", x"F7F2", x"FC9F", x"0179", x"051A", x"05B6", x"056F", x"060D", x"05F5", x"04E2", x"0431", x"0359", x"01D9", x"011A", x"0142", x"0169", x"01F6", x"02F4", x"02F4", x"01F2", x"008D", x"FEAB", x"FCF4", x"FC26", x"FB8A", x"FABF", x"FA5A", x"FA38", x"FA72", x"FBB7", x"FD93", x"FF0A", x"0046", x"00E0", x"002D", x"FF22", x"FE83", x"FDE0", x"FDB0", x"FE6C", x"FE8F", x"FD5E", x"FBB5", x"F97D", x"F6A6", x"F547", x"F5D3", x"F729", x"F91E", x"FBA7", x"FD40", x"FDE4", x"FED8", x"FF7A", x"FF48", x"FEFA", x"FE4C", x"FCBE", x"FB5F", x"FAC2", x"F9C2", x"F86E", x"F774", x"F658", x"F560", x"F59E", x"F67C", x"F6FB", x"F725", x"F719", x"F6A9", x"F617", x"F5AF", x"F55A", x"F554", x"F5B2", x"F699", x"F817", x"F96F", x"F9E8", x"FA32", x"FAAA", x"FA7B", x"F9EF", x"F9E8", x"F988", x"F885", x"F7F4", x"F75F", x"F527", x"F2B0", x"F1D5", x"F24E", x"F42E", x"F7E9", x"FBBC", x"FDC6", x"FEF3", x"FFF2", x"FFCF", x"FEB0", x"FD8D", x"FC1A", x"FA49", x"F935", x"F8E3", x"F836", x"F725", x"F683", x"F617", x"F590", x"F51B", x"F485", x"F31B", x"F156", x"F06E", x"F046", x"F014", x"EF96", x"EEE4", x"ED84", x"EC68", x"ECD2", x"EE60", x"EFB9", x"F070", x"F042", x"EEB4", x"ECA6", x"EBA0", x"EC18", x"EDC4", x"F035", x"F246", x"F251", x"F01C", x"ECE5", x"EA77", x"E9E4", x"EB5B", x"EE2C", x"F13F", x"F390", x"F509", x"F5CF", x"F586", x"F3C1", x"F16E", x"EF49", x"EDD3", x"ED93", x"EEBC", x"F061", x"F22D", x"F3DA", x"F48F", x"F391", x"F148", x"EE03", x"EA9A", x"E8AB", x"E873", x"E8E1", x"E963", x"E990", x"E8B4", x"E776", x"E78A", x"E8D3", x"EA9F", x"ECAD", x"EE52", x"EE9A", x"EDF3", x"ECE7", x"EBC1", x"EAE3", x"EAB3", x"EB1E", x"EBE5", x"EBFB", x"EA6F", x"E864", x"E722", x"E661", x"E6B2", x"E89C", x"EA74", x"EB84", x"EE2B", x"F233", x"F508", x"F6BC", x"F7F1", x"F70E", x"F4E8", x"F471", x"F515", x"F51A", x"F5CA", x"F761", x"F7DC", x"F756", x"F6E5", x"F598", x"F3AF", x"F289", x"F19F", x"EFC2", x"ED3E", x"EA5F", x"E7CD", x"E743", x"E90C", x"EBFE", x"EF4F", x"F197", x"F149", x"EF18", x"ECB2", x"EA63", x"E968", x"EA81", x"EBAC", x"EAEC", x"E88D", x"E4C0", x"E036", x"DDCB", x"DE7F", x"E05F", x"E283", x"E4A3", x"E546", x"E512", x"E630", x"E832", x"E999", x"EAF2", x"EBDD", x"EB41", x"EA63", x"EAD1", x"EB6A", x"EBC2", x"ECB5", x"EDB9", x"ED8D", x"ECE5", x"EC03", x"EA72", x"E8C4", x"E874", x"E93E", x"EA12", x"EA6A", x"EA3F", x"E9AE", x"E931", x"E9C0", x"EB9A", x"EDDD", x"EFC8", x"F176", x"F27B", x"F1EA", x"F062", x"EF44", x"EEA5", x"EE8D", x"EF81", x"F01C", x"EF14", x"ED59", x"EC77", x"EC9B", x"EE22", x"F120", x"F3CD", x"F4DB", x"F515", x"F502", x"F4B2", x"F544", x"F711", x"F908", x"FABD", x"FC7A", x"FD9E", x"FDA9", x"FD2D", x"FC4D", x"FAF9", x"F981", x"F862", x"F793", x"F72E", x"F767", x"F854", x"F9BB", x"FA66", x"F9DD", x"F8E5", x"F7EC", x"F6A8", x"F616", x"F6B1", x"F6F4", x"F6C0", x"F759", x"F778", x"F53F", x"F29A", x"F177", x"F130", x"F25B", x"F5A7", x"F7C7", x"F65A", x"F417", x"F302", x"F2C3", x"F458", x"F811", x"FA91", x"FAA2", x"FA5E", x"FA0D", x"F90D", x"F8C8", x"F914", x"F837", x"F711", x"F715", x"F774", x"F7BD", x"F8A3", x"F8F4", x"F7DE", x"F69D", x"F578", x"F380", x"F16D", x"F014", x"EF1C", x"EE8E", x"EE59", x"EDC7", x"ECE2", x"EC44", x"EC12", x"ECDA", x"EE5C", x"EF03", x"EEB5", x"EE73", x"ECC4", x"E98A", x"E794", x"E7B5", x"E866", x"EAD2", x"EE42", x"EE5B", x"EAE6", x"E801", x"E625", x"E4F2", x"E6CD", x"EA8F", x"EC3D", x"ECCF", x"EE4C", x"EF0D", x"EF47", x"F114", x"F30B", x"F3A0", x"F497", x"F5AA", x"F579", x"F567", x"F62D", x"F642", x"F613", x"F65C", x"F5A3", x"F430", x"F3AE", x"F3B2", x"F419", x"F5DE", x"F771", x"F775", x"F71D", x"F677", x"F533", x"F593", x"F7C1", x"F97C", x"FB1B", x"FD06", x"FC7A", x"FA5E", x"FA40", x"FB60", x"FC86", x"FF3F", x"015F", x"FEFF", x"FACD", x"F87E", x"F736", x"F7FA", x"FC1E", x"FF95", x"FF99", x"FEBF", x"FE04", x"FCC8", x"FD76", x"0049", x"0212", x"02E2", x"043B", x"04BF", x"04E6", x"0671", x"07B3", x"0754", x"0729", x"070D", x"05CD", x"050E", x"0550", x"04E9", x"04B8", x"061A", x"0773", x"0878", x"0A39", x"0B3D", x"0B0C", x"0B65", x"0C2F", x"0C6A", x"0D90", x"0F44", x"0F33", x"0E57", x"0E45", x"0DBD", x"0CA7", x"0C49", x"0AA3", x"0622", x"01B7", x"FF4D", x"FE4A", x"FF17", x"01F2", x"03FB", x"043E", x"042E", x"043C", x"03EF", x"042E", x"0562", x"06BE", x"07D2", x"08B7", x"08E7", x"0888", x"07FF", x"079F", x"0740", x"0666", x"04D6", x"0319", x"01DF", x"016F", x"0215", x"0362", x"0400", x"03DC", x"03BD", x"0391", x"0351", x"03CA", x"045C", x"03E6", x"033B", x"0329", x"0257", x"007E", x"FF18", x"FE45", x"FD8A", x"FDF6", x"FF87", x"FFE3", x"FEA5", x"FE07", x"FEA1", x"FFEE", x"0232", x"054F", x"0752", x"07D3", x"07C5", x"0712", x"0519", x"02DE", x"01CA", x"01FF", x"02EC", x"046C", x"061A", x"0795", x"092C", x"0B53", x"0D7D", x"0E73", x"0DDC", x"0C21", x"09E2", x"07E7", x"0744", x"07F0", x"08F2", x"09F8", x"0AC3", x"0ADC", x"0ABB", x"0BB4", x"0CF1", x"0D88", x"0E63", x"0F6B", x"0EBC", x"0D4B", x"0CAE", x"0BDA", x"0ADA", x"0C49", x"0E83", x"0DA3", x"0B12", x"098B", x"082E", x"0823", x"0B88", x"0EEB", x"0E87", x"0CE7", x"0C0E", x"0A77", x"097C", x"0AD0", x"0BF9", x"0C36", x"0DC9", x"0FC6", x"102B", x"1042", x"1068", x"0F58", x"0EA9", x"0F8D", x"103F", x"10AA", x"11BC", x"11F5", x"1120", x"1158", x"1260", x"12BA", x"1315", x"1318", x"1145", x"0F68", x"0F1F", x"0F5F", x"0FE3", x"10CD", x"1052", x"0E75", x"0D9A", x"0DF0", x"0F2A", x"1245", x"1539", x"14D4", x"1234", x"0F59", x"0C2D", x"0AD9", x"0CF8", x"0F1A", x"0EA1", x"0D3D", x"0B07", x"078C", x"05D1", x"06FC", x"0877", x"09EA", x"0C55", x"0D9F", x"0D35", x"0D5F", x"0E2D", x"0E81", x"0F7D", x"10C7", x"104C", x"0EA2", x"0D31", x"0BAC", x"0AEA", x"0C29", x"0E19", x"0F90", x"10CA", x"1163", x"1142", x"1204", x"13E4", x"1578", x"16A9", x"1714", x"15A7", x"13B9", x"1307", x"12FE", x"130D", x"1390", x"12BF", x"0F81", x"0C09", x"09D0", x"08A7", x"09AD", x"0D4E", x"10CE", x"132F", x"158B", x"173B", x"1749", x"1752", x"179C", x"16DD", x"1608", x"1652", x"1625", x"14E7", x"13C3", x"129B", x"10E4", x"0FCD", x"0FA3", x"0EBD", x"0D2C", x"0C4A", x"0C3A", x"0CE6", x"0E88", x"1071", x"1172", x"11BE", x"1225", x"12E5", x"13A0", x"1391", x"1283", x"107E", x"0DB6", x"0ABA", x"08D0", x"0831", x"083D", x"0913", x"0A84", x"0B3E", x"0B10", x"0B9C", x"0D27", x"0EBE", x"1088", x"1208", x"1201", x"10AB", x"0F57", x"0DF5", x"0C43", x"0ADE", x"09FF", x"0943", x"08C2", x"0888", x"087D", x"08F7", x"0A38", x"0BC3", x"0D27", x"0DA9", x"0CB9", x"0AC9", x"08B2", x"068C", x"050B", x"04DA", x"0580", x"0681", x"07A5", x"07FF", x"0707", x"0603", x"05AC", x"05C8", x"073B", x"099E", x"0AD1", x"0A91", x"0A40", x"096F", x"086D", x"0912", x"0A1F", x"08CB", x"0626", x"03FF", x"01CF", x"0113", x"03A8", x"06E5", x"0842", x"092B", x"0A0D", x"09AE", x"09C2", x"0BAD", x"0D42", x"0DEB", x"0F04", x"0F80", x"0E2F", x"0CC3", x"0C0A", x"0B52", x"0B2D", x"0C03", x"0C53", x"0B91", x"0AAE", x"09F8", x"09A3", x"0A04", x"0AB0", x"0B44", x"0BE4", x"0C6A", x"0D19", x"0E5E", x"0FA8", x"107A", x"11A6", x"12C6", x"12AE", x"120B", x"119A", x"10D8", x"1013", x"106E", x"10A7", x"0FBA", x"0ECE", x"0EB3", x"0ECB", x"0F7D", x"10E2", x"1189", x"110E", x"1039", x"0F6B", x"0E8D", x"0E6C", x"0F48", x"10D3", x"12F1", x"156A", x"17D8", x"19F8", x"1BBF", x"1D7C", x"1F12", x"1FB7", x"1EF8", x"1CFC", x"19B0", x"15D3", x"136E", x"12EA", x"12E7", x"1370", x"14D1", x"157A", x"153A", x"15D7", x"16B2", x"1696", x"179C", x"1ACE", x"1D99", x"1EEC", x"200C", x"1FF9", x"1E67", x"1D8F", x"1DDA", x"1C87", x"19C7", x"17B2", x"16B3", x"1692", x"181C", x"1A5B", x"1B84", x"1BBA", x"1C03", x"1C40", x"1C5C", x"1CAD", x"1D30", x"1D96", x"1DBB", x"1DB0", x"1D63", x"1CFF", x"1C74", x"1B8F", x"19E9", x"1760", x"146F", x"11A1", x"0F75", x"0E75", x"0EC1", x"0F7A", x"1008", x"1064", x"1038", x"0F78", x"0F1F", x"0F9E", x"0FD9", x"0F77", x"0F6E", x"0FAD", x"0F7E", x"0F3A", x"0F14", x"0E45", x"0CE1", x"0C5D", x"0CAF", x"0C7F", x"0C02", x"0C49", x"0D06", x"0DE7", x"0F3A", x"10C7", x"113D", x"106F", x"0EBB", x"0C02", x"0868", x"0531", x"0392", x"03BC", x"0522", x"06E7", x"08C6", x"0AA7", x"0C2E", x"0D51", x"0E97", x"0F87", x"0F76", x"0F1E", x"0EB3", x"0D2F", x"0B0D", x"09C3", x"08E6", x"07D0", x"073F", x"0692", x"04C2", x"0300", x"0266", x"021E", x"02E1", x"054A", x"071F", x"0771", x"081C", x"0883", x"07AC", x"075D", x"0747", x"04A4", x"019B", x"01AE", x"032D", x"0482", x"06C7", x"07BE", x"052C", x"02C7", x"0321", x"035C", x"0325", x"03C4", x"031E", x"008D", x"FF4F", x"FF91", x"FF35", x"FF48", x"0027", x"FFB3", x"FEC6", x"FF18", x"FFBA", x"FFEC", x"00AF", x"0134", x"00A2", x"0061", x"00A7", x"006D", x"0010", x"FFAF", x"FEB4", x"FDBB", x"FD00", x"FBDE", x"FAEC", x"FA7C", x"F923", x"F781", x"F724", x"F706", x"F6AB", x"F7B4", x"F88F", x"F707", x"F5BB", x"F6A9", x"F790", x"F864", x"FAB1", x"FC4B", x"FB98", x"FB72", x"FBD6", x"FA3E", x"F7F5", x"F75C", x"F7A5", x"F875", x"FAEF", x"FD8C", x"FEBB", x"FF76", x"0045", x"0095", x"0096", x"0085", x"FFDD", x"FE90", x"FCA5", x"FA00", x"F779", x"F5C8", x"F4F2", x"F56F", x"F6F3", x"F825", x"F8FC", x"F9E8", x"F9D9", x"F923", x"F980", x"FA26", x"FA23", x"FB39", x"FD31", x"FDA4", x"FD4A", x"FD31", x"FAD1", x"F6D6", x"F5CA", x"F7C2", x"FA3B", x"FE04", x"0224", x"0307", x"01FA", x"02BE", x"03BF", x"0325", x"02BF", x"0257", x"0055", x"FED2", x"FF1F", x"FEF7", x"FDE9", x"FD42", x"FC18", x"FA2D", x"F91A", x"F887", x"F761", x"F6AC", x"F66E", x"F5F7", x"F666", x"F849", x"FA1A", x"FB64", x"FC95", x"FC88", x"FB34", x"FA0C", x"F89A", x"F656", x"F47D", x"F36A", x"F24B", x"F24C", x"F383", x"F3F7", x"F35F", x"F2A2", x"F0EF", x"EF0D", x"EFEA", x"F305", x"F5FE", x"F8C1", x"FAAF", x"F9DB", x"F78E", x"F65A", x"F52E", x"F37B", x"F29D", x"F25F", x"F15A", x"F0D1", x"F187", x"F252", x"F336", x"F484", x"F4C5", x"F34E", x"F12E", x"EEC6", x"EC66", x"EAE0", x"E9EB", x"E8B5", x"E7B9", x"E71C", x"E68D", x"E677", x"E70C", x"E786", x"E7F1", x"E860", x"E852", x"E830", x"E8CA", x"E955", x"E998", x"EA32", x"EA36", x"E8F3", x"E7A0", x"E5DF", x"E29C", x"DFDB", x"DFBF", x"E0D9", x"E298", x"E58D", x"E79B", x"E798", x"E822", x"EA26", x"EB3C", x"EBC5", x"ECC4", x"ED1D", x"ECE6", x"EE34", x"EFED", x"F021", x"EF9C", x"EEF0", x"ED89", x"EC41", x"EC03", x"EB9E", x"EAFF", x"EADA", x"EB1D", x"EBD7", x"ED5D", x"EEF3", x"EFF9", x"F0D6", x"F12B", x"F107", x"F152", x"F1A1", x"F16C", x"F1F4", x"F33E", x"F3AE", x"F43F", x"F5F8", x"F6B9", x"F617", x"F5A4", x"F3FA", x"F03E", x"EEBF", x"F116", x"F414", x"F6C2", x"F97F", x"F933", x"F60B", x"F4CE", x"F5FA", x"F637", x"F648", x"F721", x"F6D5", x"F636", x"F7F6", x"FABE", x"FC31", x"FD51", x"FE4A", x"FD95", x"FBD8", x"FA53", x"F89A", x"F6E6", x"F626", x"F5F4", x"F566", x"F44C", x"F29E", x"F0D1", x"EFF5", x"F081", x"F280", x"F5A6", x"F8C2", x"FB31", x"FD6C", x"FEFC", x"FF6D", x"FFAD", x"FFC1", x"FE88", x"FC9A", x"FAA3", x"F744", x"F34C", x"F175", x"F1C2", x"F2E1", x"F560", x"F823", x"F878", x"F714", x"F602", x"F456", x"F210", x"F167", x"F253", x"F39C", x"F5C7", x"F851", x"F924", x"F850", x"F70E", x"F549", x"F385", x"F275", x"F18E", x"F09F", x"F045", x"EFC9", x"EED6", x"EE2C", x"ED44", x"EB98", x"EAAB", x"EAA3", x"EA1B", x"E9CA", x"EA3C", x"E999", x"E81E", x"E7B4", x"E76F", x"E6DC", x"E841", x"EB1D", x"EC93", x"ED0B", x"ECC0", x"EA02", x"E6EE", x"E765", x"EA18", x"EC8D", x"EF12", x"EFCB", x"ECDB", x"E942", x"E755", x"E526", x"E28B", x"E131", x"E001", x"DEEC", x"E04F", x"E384", x"E602", x"E83F", x"E9FD", x"E9F9", x"E94F", x"E99A", x"E9D6", x"EA12", x"EB2D", x"EBE2", x"EB80", x"EB84", x"EB86", x"EA73", x"E937", x"E804", x"E5EF", x"E43D", x"E444", x"E51F", x"E6B8", x"E99D", x"EC81", x"EEE1", x"F1A5", x"F3D3", x"F41C", x"F319", x"F0F5", x"ED81", x"EB4C", x"EBF9", x"EE0B", x"F079", x"F305", x"F3D8", x"F2C9", x"F212", x"F253", x"F2C3", x"F3EA", x"F5AE", x"F6E3", x"F741", x"F753", x"F6DC", x"F6CB", x"F79F", x"F8AA", x"F94E", x"F8E2", x"F650", x"F306", x"F165", x"F0ED", x"F105", x"F293", x"F41D", x"F3D3", x"F3DE", x"F4F7", x"F498", x"F38B", x"F43E", x"F4D3", x"F4AA", x"F65B", x"F859", x"F80D", x"F862", x"FB02", x"FC96", x"FCA6", x"FCA5", x"F982", x"F38A", x"F0AF", x"F1E1", x"F3D2", x"F6A0", x"F96A", x"F819", x"F409", x"F1C4", x"F043", x"EDFE", x"ED0E", x"ED0F", x"EBDC", x"EB4B", x"EC9F", x"ED92", x"EE28", x"EFC2", x"F132", x"F196", x"F218", x"F1D6", x"F059", x"EF6F", x"EF5F", x"EF64", x"F07B", x"F2AA", x"F3BC", x"F433", x"F4C7", x"F431", x"F2BA", x"F2BD", x"F33E", x"F30D", x"F38C", x"F4E3", x"F590", x"F6D6", x"F958", x"FA37", x"F892", x"F5F3", x"F24A", x"EEC3", x"EEC6", x"F232", x"F65A", x"FA81", x"FDDF", x"FE41", x"FCCE", x"FBE7", x"FB00", x"FA1C", x"FACE", x"FC89", x"FDC5", x"FF1E", x"0052", x"0011", x"FF05", x"FE2E", x"FCBE", x"FAD5", x"F943", x"F79E", x"F668", x"F6A3", x"F72C", x"F76C", x"F821", x"F89E", x"F835", x"F838", x"F85C", x"F6F8", x"F5DC", x"F677", x"F706", x"F73A", x"F82A", x"F7CD", x"F5BE", x"F57D", x"F73A", x"F85D", x"F9B1", x"FB0D", x"F9EA", x"F80F", x"F8E6", x"FAB8", x"FBDF", x"FDAD", x"FE56", x"FBDA", x"F947", x"F838", x"F672", x"F4C1", x"F49B", x"F3D8", x"F285", x"F326", x"F4A5", x"F533", x"F688", x"F839", x"F898", x"F94E", x"FAF3", x"FB22", x"FA6D", x"FA53", x"F972", x"F843", x"F920", x"FA24", x"F955", x"F860", x"F70E", x"F40F", x"F214", x"F278", x"F25B", x"F1CB", x"F27A", x"F334", x"F41B", x"F7BA", x"FC44", x"FE73", x"FEED", x"FDE7", x"FAEB", x"F931", x"FB11", x"FE7F", x"023E", x"05FB", x"070F", x"050D", x"0302", x"018B", x"0059", x"013B", x"0395", x"0501", x"0630", x"07CE", x"0803", x"0758", x"073C", x"0622", x"03E9", x"029F", x"019E", x"FFC2", x"FEF0", x"FEFD", x"FE27", x"FDF6", x"FF73", x"004F", x"008E", x"01C5", x"023F", x"01CD", x"0308", x"055C", x"0687", x"07D7", x"09A1", x"0A59", x"0B62", x"0E52", x"1090", x"10A5", x"0FF1", x"0E20", x"0B7F", x"0B1B", x"0D58", x"0F7A", x"10DA", x"1158", x"0F44", x"0BB3", x"093A", x"07D9", x"070E", x"07F6", x"0A03", x"0BBC", x"0DA6", x"0FC2", x"1139", x"124A", x"13D2", x"152D", x"1620", x"16B9", x"1639", x"149C", x"12DE", x"113C", x"101B", x"1058", x"1179", x"1234", x"12BA", x"12C8", x"11D0", x"1124", x"1201", x"134C", x"1473", x"15BE", x"166C", x"163B", x"1710", x"18E0", x"19F8", x"1A1A", x"1981", x"1766", x"1535", x"155E", x"177D", x"1A26", x"1D4F", x"1F68", x"1EC6", x"1CB9", x"1B05", x"193C", x"17E5", x"180E", x"1897", x"187C", x"18C8", x"1938", x"18BA", x"17FE", x"17B8", x"16D9", x"1595", x"14A5", x"134D", x"119C", x"110C", x"1187", x"1270", x"1443", x"1640", x"16AD", x"15EA", x"14D8", x"12E0", x"10D4", x"1026", x"0FAB", x"0E88", x"0DBF", x"0DA4", x"0D5F", x"0DEE", x"0F3C", x"0F77", x"0E5C", x"0D4F", x"0C96", x"0CCD", x"0F33", x"12EB", x"163C", x"18A3", x"193C", x"1753", x"142A", x"111C", x"0E3A", x"0C5F", x"0C2C", x"0C35", x"0C58", x"0D5F", x"0E7F", x"0F15", x"1023", x"1169", x"11C4", x"1240", x"1355", x"13B9", x"13C6", x"14A0", x"1537", x"155F", x"1647", x"16D4", x"15A6", x"13C1", x"11A0", x"0ECE", x"0CDD", x"0CDE", x"0CEA", x"0C92", x"0CF2", x"0D85", x"0E41", x"1049", x"1283", x"12E2", x"1215", x"1121", x"102A", x"10C0", x"13C4", x"1757", x"1A83", x"1D42", x"1E0B", x"1C95", x"1A77", x"17C9", x"1430", x"11AE", x"10E7", x"1092", x"11A8", x"1479", x"166F", x"169E", x"167F", x"1557", x"1303", x"11F5", x"122A", x"1190", x"1103", x"1163", x"1108", x"100E", x"0FC6", x"0E5F", x"0AF7", x"080F", x"0680", x"0585", x"0666", x"08B5", x"0971", x"0875", x"07D7", x"0751", x"06CF", x"0788", x"0822", x"069E", x"0470", x"0347", x"02DD", x"03C1", x"0688", x"0978", x"0B20", x"0BD7", x"0B5A", x"0954", x"0724", x"05F8", x"05EF", x"070D", x"08BC", x"09DF", x"09FF", x"097A", x"08C3", x"08C7", x"09C8", x"0B28", x"0C9B", x"0DBD", x"0D8E", x"0C0E", x"0A30", x"07EB", x"05B3", x"0536", x"0668", x"07EA", x"09B8", x"0B4E", x"0B24", x"09C8", x"0926", x"08D8", x"089F", x"09C0", x"0B9E", x"0D01", x"0E7F", x"1043", x"10A7", x"0FE1", x"0F28", x"0E0F", x"0CF5", x"0D76", x"0ECA", x"0FD9", x"10F4", x"116E", x"1018", x"0E80", x"0DEA", x"0DA1", x"0E0B", x"0FFF", x"11B2", x"1277", x"13BF", x"14FC", x"14FC", x"14FA", x"1581", x"14FF", x"1402", x"1373", x"1237", x"1065", x"0FAF", x"0FC6", x"0FCC", x"105D", x"10E8", x"1038", x"0F36", x"0E89", x"0D76", x"0C8E", x"0C67", x"0BC3", x"0A8A", x"0A02", x"0A08", x"0A1B", x"0B03", x"0BD0", x"0B37", x"0A10", x"09AF", x"0A10", x"0BF9", x"0F7C", x"12F8", x"157B", x"16F7", x"1695", x"146C", x"124B", x"103C", x"0E82", x"0E1A", x"0E6B", x"0DDD", x"0D73", x"0DAF", x"0D11", x"0BFB", x"0B95", x"0ABF", x"099E", x"0A79", x"0C7C", x"0DA0", x"0E9B", x"0F61", x"0E44", x"0CE7", x"0D0A", x"0CE2", x"0B9A", x"0AF9", x"0A0D", x"07FC", x"072B", x"07A7", x"069C", x"0499", x"037D", x"0269", x"01D3", x"03DC", x"0691", x"0709", x"0627", x"0508", x"030E", x"0191", x"0256", x"03C8", x"0480", x"04F2", x"0470", x"0218", x"FF0F", x"FCC5", x"FB7A", x"FBA8", x"FD5D", x"FF9B", x"01AC", x"03B2", x"0553", x"06C7", x"084B", x"0969", x"09F6", x"0A67", x"0A4F", x"0930", x"07E4", x"06CA", x"0589", x"04B8", x"048E", x"0379", x"00DF", x"FDEE", x"FB25", x"F8DB", x"F898", x"FA9E", x"FD17", x"FF88", x"027C", x"04CE", x"0598", x"05C0", x"0556", x"0401", x"034B", x"04C8", x"0770", x"0A47", x"0D58", x"0FAE", x"104A", x"0FD4", x"0E99", x"0C0B", x"0881", x"0556", x"02EF", x"0175", x"014E", x"020D", x"02DE", x"038D", x"0430", x"04BB", x"0573", x"0685", x"0829", x"0A47", x"0C6E", x"0E1A", x"0F13", x"0ED9", x"0D52", x"0BA3", x"0A43", x"08C7", x"0796", x"0735", x"06B8", x"0605", x"0653", x"06AC", x"05C8", x"0503", x"0557", x"057E", x"059B", x"0673", x"065D", x"04CA", x"0463", x"05BA", x"0735", x"08EC", x"0ADF", x"0B2C", x"09E9", x"08C4", x"074B", x"050D", x"0382", x"02DF", x"026B", x"02B2", x"0382", x"03BC", x"03BC", x"0416", x"040D", x"03E3", x"047D", x"050A", x"0523", x"057D", x"054A", x"03BE", x"0237", x"013D", x"0012", x"FF7E", x"FF7E", x"FE59", x"FC0B", x"F9FA", x"F7DF", x"F5C5", x"F550", x"F55F", x"F46D", x"F3BE", x"F437", x"F443", x"F425", x"F495", x"F3EC", x"F236", x"F241", x"F490", x"F778", x"FB16", x"FF21", x"018E", x"020E", x"01AA", x"0028", x"FD61", x"FAC5", x"F92F", x"F808", x"F6AD", x"F4B4", x"F277", x"F099", x"EF81", x"EF64", x"F039", x"F0CF", x"F0D2", x"F1A9", x"F342", x"F460", x"F552", x"F6E8", x"F7FC", x"F8E9", x"FB09", x"FCE8", x"FCA9", x"FBE6", x"FB6E", x"FA17", x"F8AA", x"F81B", x"F65B", x"F30E", x"F0D4", x"EFB5", x"EE39", x"ED49", x"ED46", x"ECA5", x"ECB7", x"EF9D", x"F3D2", x"F778", x"FAC4", x"FCE0", x"FCB8", x"FBEF", x"FBA2", x"FB0F", x"FA74", x"FAC8", x"FB3E", x"FB7E", x"FC0D", x"FC68", x"FC32", x"FC2F", x"FC25", x"FB81", x"FB4D", x"FB92", x"FBD6", x"FC93", x"FD84", x"FCF5", x"FB4B", x"FA37", x"F926", x"F803", x"F7E4", x"F74B", x"F4E4", x"F326", x"F37F", x"F41F", x"F51E", x"F6EE", x"F705", x"F583", x"F5DB", x"F7D1", x"F896", x"F8EA", x"F8EB", x"F6C0", x"F455", x"F498", x"F5D4", x"F656", x"F781", x"F882", x"F7AA", x"F622", x"F47E", x"F189", x"EE6E", x"ED06", x"EC7B", x"EC81", x"ED3C", x"ED29", x"EBA9", x"EA13", x"E828", x"E5E2", x"E53C", x"E615", x"E6D2", x"E809", x"E9A3", x"E9CB", x"E986", x"EAA8", x"EB93", x"EB4F", x"EB48", x"EA66", x"E7D8", x"E6B3", x"E7B0", x"E87F", x"E95A", x"EA83", x"E95B", x"E6B0", x"E609", x"E641", x"E595", x"E5D2", x"E689", x"E5ED", x"E68E", x"EA10", x"ED29", x"EEB1", x"F02C", x"F04B", x"EE89", x"ED60", x"ED11", x"EC16", x"EBA7", x"ECCC", x"EE07", x"EF65", x"F131", x"F24F", x"F2A1", x"F2D5", x"F1ED", x"EFD4", x"EE08", x"EC35", x"EA1F", x"E90C", x"E82E", x"E642", x"E501", x"E56B", x"E5DC", x"E68F", x"E7F9", x"E7F3", x"E647", x"E55D", x"E4F8", x"E435", x"E4E0", x"E6DD", x"E83F", x"E9F4", x"EC6E", x"ECEB", x"EAE5", x"E80F", x"E431", x"E025", x"DF5A", x"E1BB", x"E4C1", x"E84C", x"EBC5", x"ED0F", x"ECAF", x"EC6B", x"EB39", x"E8FC", x"E760", x"E639", x"E4DF", x"E478", x"E4A3", x"E415", x"E328", x"E203", x"DFEE", x"DE1A", x"DDD5", x"DE69", x"DFDA", x"E22A", x"E35A", x"E2E1", x"E296", x"E24F", x"E177", x"E14B", x"E12E", x"DF4E", x"DD5D", x"DD43", x"DD80", x"DDFB", x"DFDE", x"E10A", x"E075", x"E0DC", x"E26A", x"E305", x"E3DD", x"E5B5", x"E6A1", x"E764", x"EA2B", x"ED2A", x"EE8A", x"EFB4", x"F009", x"EE53", x"EC8A", x"EBE6", x"EA98", x"E925", x"E8CE", x"E81A", x"E70C", x"E752", x"E7E4", x"E783", x"E7A7", x"E87A", x"E90F", x"EACE", x"EDED", x"F00A", x"F09A", x"F0AB", x"EF6D", x"ED7E", x"ED14", x"ED48", x"ECF7", x"ECF6", x"ECCD", x"EB32", x"EA10", x"EA45", x"EA0C", x"E9D8", x"EA8D", x"EA41", x"E93E", x"EA8A", x"ECFB", x"EE20", x"EF3C", x"F031", x"EF5D", x"EF6B", x"F2DD", x"F6B9", x"F925", x"FB49", x"FBB4", x"F952", x"F719", x"F589", x"F29C", x"EF69", x"EDA9", x"EC21", x"EB8C", x"ED49", x"EFA0", x"F13F", x"F326", x"F4A5", x"F4E5", x"F5D5", x"F799", x"F8E8", x"FAB6", x"FD68", x"FF13", x"001B", x"017E", x"017B", x"FFFA", x"FEFA", x"FDAE", x"FBA3", x"FB47", x"FC38", x"FC1C", x"FC34", x"FCC5", x"FB70", x"F9BA", x"FA2D", x"FA55", x"F8EA", x"F8BE", x"F99E", x"FAB4", x"FF88", x"0814", x"0ED9", x"1251", x"13F0", x"123F", x"0E47", x"0C5D", x"0BF8", x"0A86", x"098D", x"09F1", x"09D8", x"09DF", x"0B41", x"0BD6", x"0B18", x"0A45", x"08FD", x"0700", x"05EA", x"05C0", x"05FB", x"0732", x"0886", x"08A2", x"08E2", x"09B6", x"0A04", x"0A83", x"0B43", x"09E9", x"070C", x"0552", x"03BA", x"01A6", x"0121", x"0146", x"FFF5", x"FF67", x"0025", x"FEEE", x"FBF3", x"F9D4", x"F7CF", x"F6B5", x"F9EC", x"FFE0", x"04E2", x"094B", x"0D28", x"0E42", x"0E34", x"0EEC", x"0E96", x"0CCB", x"0BB3", x"0A8E", x"088C", x"0769", x"0696", x"042B", x"0169", x"FF1C", x"FC25", x"F9E6", x"F9A4", x"F98A", x"F94B", x"FA47", x"FB26", x"FBA2", x"FDE5", x"00F9", x"0274", x"035D", x"03EC", x"0267", x"00FA", x"01DF", x"028D", x"01D8", x"01A4", x"00C6", x"FE5A", x"FD9A", x"FE7A", x"FDCE", x"FC71", x"FC78", x"FCDC", x"FE7D", x"0378", x"0926", x"0C5C", x"0DED", x"0DCB", x"0B3F", x"08D9", x"082F", x"07CD", x"07CC", x"089A", x"0890", x"0782", x"0700", x"064E", x"04F2", x"0453", x"03F5", x"02F0", x"02FF", x"0465", x"0554", x"0660", x"07FA", x"083F", x"0777", x"075D", x"069E", x"047B", x"02EF", x"017E", x"FF18", x"FD9A", x"FD78", x"FC62", x"FB04", x"FAC0", x"FA12", x"F956", x"FA95", x"FBCB", x"FACB", x"F935", x"F791", x"F58F", x"F616", x"FA4B", x"FECB", x"0212", x"0460", x"0421", x"01BC", x"0098", x"0098", x"0021", x"0039", x"00AF", x"FF97", x"FE42", x"FDD7", x"FC6B", x"F9F3", x"F813", x"F5EF", x"F36E", x"F2B3", x"F358", x"F3A7", x"F4DA", x"F716", x"F8A6", x"FA70", x"FD50", x"FF42", x"FFF6", x"00DB", x"010B", x"0068", x"0148", x"035F", x"04DB", x"069F", x"0890", x"08DD", x"084B", x"087C", x"07B0", x"05E3", x"055D", x"05FF", x"075E", x"0B21", x"105F", x"13FD", x"15D1", x"16A7", x"1567", x"1316", x"11A7", x"1038", x"0E24", x"0D1E", x"0D5D", x"0E22", x"1010", x"1298", x"1398", x"12EA", x"1146", x"0E70", x"0B7D", x"0996", x"0861", x"0793", x"07D4", x"0837", x"0857", x"0957", x"0AA3", x"0B10", x"0B49", x"0B18", x"0923", x"06E0", x"0634", x"05FC", x"0604", x"07C4", x"09BD", x"0A7C", x"0B5C", x"0C31", x"0A88", x"07AF", x"05D7", x"04B5", x"050C", x"0896", x"0D31", x"100C", x"11C4", x"1296", x"11BA", x"10EB", x"116A", x"1165", x"103A", x"0EFA", x"0CF8", x"0A25", x"083A", x"072A", x"05DB", x"04F9", x"04A5", x"03C1", x"02EC", x"030A", x"030F", x"0366", x"04DD", x"0697", x"07E2", x"09D7", x"0B95", x"0BA5", x"0B44", x"0AEA", x"09C3", x"08ED", x"09CB", x"0A50", x"09B1", x"0975", x"095B", x"087F", x"083B", x"0865", x"06C1", x"0416", x"02A3", x"028B", x"03F6", x"07B5", x"0BB6", x"0D81", x"0D7F", x"0C5D", x"0A63", x"092D", x"09B8", x"0A85", x"0AEA", x"0B22", x"0ABB", x"0A2A", x"0AEB", x"0C90", x"0E30", x"0FB7", x"10AB", x"105C", x"1007", x"107B", x"1137", x"128E", x"144F", x"14D2", x"13E3", x"1283", x"1015", x"0CAF", x"09ED", x"077C", x"0490", x"02C6", x"026B", x"01C0", x"016A", x"02E7", x"04B0", x"0637", x"089F", x"0A1D", x"0923", x"0838", x"0905", x"0AE5", x"0E83", x"13F4", x"17D8", x"1917", x"1996", x"1921", x"17DB", x"17B0", x"1826", x"16E0", x"14AE", x"1264", x"0F12", x"0BBB", x"0A0D", x"0843", x"05A9", x"03E6", x"02FC", x"0265", x"03E1", x"074D", x"0A5D", x"0D3B", x"1045", x"124B", x"13A8", x"15F6", x"17DC", x"1896", x"1938", x"1916", x"175A", x"15DC", x"1523", x"13CE", x"1301", x"13B6", x"1426", x"13A2", x"130F", x"10FA", x"0D16", x"0A80", x"0ABC", x"0CFE", x"11A6", x"17AF", x"1BF0", x"1DAA", x"1E1C", x"1D3D", x"1B8C", x"1AAC", x"1A40", x"196F", x"18E5", x"18B8", x"1826", x"17EE", x"1802", x"1758", x"166E", x"15AD", x"148A", x"13A4", x"13E5", x"1412", x"13EE", x"147B", x"14D0", x"1464", x"150E", x"1653", x"1639", x"158C", x"14F6", x"12AC", x"0FBB", x"0E73", x"0D39", x"0B24", x"0A8D", x"0B64", x"0BAD", x"0CB4", x"0E47", x"0D5D", x"0A87", x"08E3", x"0850", x"093F", x"0D70", x"12CE", x"15F6", x"179C", x"1833", x"16D9", x"159C", x"162B", x"161E", x"14D6", x"13B5", x"11D3", x"0EC0", x"0CC1", x"0B71", x"08D3", x"0663", x"053B", x"0416", x"03F1", x"060F", x"0865", x"0A11", x"0C83", x"0EB7", x"0FB3", x"1146", x"12F7", x"127D", x"10FA", x"0F89", x"0D10", x"0ACF", x"0B0B", x"0BC2", x"0B8B", x"0C52", x"0D7C", x"0D0B", x"0C0D", x"0AC8", x"0764", x"0360", x"0230", x"03A1", x"06E4", x"0C2B", x"114A", x"13F2", x"150A", x"15C3", x"15EF", x"16C0", x"18C5", x"1A65", x"1B53", x"1C05", x"1C01", x"1B70", x"1B69", x"1B2B", x"19F1", x"1892", x"174D", x"15C4", x"1540", x"15FB", x"16EC", x"17DE", x"18CE", x"1858", x"16E5", x"15A7", x"144C", x"12CB", x"121C", x"114E", x"0F92", x"0E69", x"0E24", x"0D5D", x"0D1A", x"0E69", x"0FC0", x"1104", x"130F", x"13FC", x"1293", x"1103", x"105A", x"1030", x"11B3", x"14C5", x"16CD", x"1761", x"17AA", x"16E7", x"1570", x"14C5", x"13B2", x"10DE", x"0D90", x"0A13", x"05D6", x"02BA", x"017E", x"FFA8", x"FD24", x"FB4B", x"F943", x"F744", x"F7AD", x"F9BD", x"FB4A", x"FD92", x"00D2", x"02EF", x"0450", x"0608", x"060B", x"0403", x"02C1", x"021B", x"010D", x"0101", x"020A", x"01D5", x"0163", x"0280", x"0337", x"0234", x"007A", x"FD8C", x"F936", x"F6BD", x"F7E8", x"FB0B", x"FF09", x"03B7", x"0705", x"087A", x"0991", x"0A91", x"0A9E", x"0A5C", x"0A18", x"093D", x"07EA", x"06BE", x"0570", x"03D3", x"026E", x"0148", x"003D", x"FF81", x"FF56", x"FFB0", x"00AF", x"021B", x"0396", x"04B2", x"04C1", x"03D7", x"027C", x"00C7", x"FEB4", x"FCBC", x"FB0B", x"F94F", x"F84A", x"F889", x"F93A", x"F9D0", x"FAA1", x"FB41", x"FAF2", x"FA13", x"F8BA", x"F668", x"F40E", x"F31A", x"F3AF", x"F59B", x"F88F", x"FB25", x"FC4B", x"FC44", x"FBA7", x"FAC8", x"FB02", x"FC28", x"FCCB", x"FC3E", x"FABC", x"F7D4", x"F45B", x"F1E9", x"EFEC", x"ED6C", x"EB38", x"E9CA", x"E886", x"E841", x"E9A3", x"EB16", x"EC20", x"EDBF", x"EF3E", x"F005", x"F115", x"F228", x"F1A9", x"F094", x"EFC4", x"EE2E", x"EC9A", x"ECAB", x"ED34", x"ED85", x"EF99", x"F2B6", x"F44D", x"F464", x"F35F", x"EFBF", x"EB92", x"EAA7", x"EC82", x"EF10", x"F288", x"F57A", x"F5E0", x"F562", x"F5D6", x"F5F8", x"F5A3", x"F5F6", x"F5CD", x"F477", x"F35C", x"F27D", x"F0F3", x"F002", x"F044", x"F08C", x"F126", x"F259", x"F296", x"F182", x"F0A4", x"EFF2", x"EF9C", x"F0B6", x"F2AC", x"F3E9", x"F498", x"F4BD", x"F37B", x"F163", x"EF4C", x"ECAB", x"EA38", x"E93A", x"E921", x"E998", x"EB8E", x"EDF0", x"EEFF", x"EF1E", x"EE79", x"EC76", x"EB2A", x"ECA4", x"EFCB", x"F324", x"F6A9", x"F8FE", x"F95F", x"F988", x"FA27", x"FA5A", x"FA10", x"F98C", x"F7D1", x"F537", x"F2A6", x"F00B", x"EDB6", x"EC68", x"EB93", x"EAE9", x"EB1E", x"EBB5", x"EC35", x"ED79", x"EF3F", x"F087", x"F209", x"F46E", x"F655", x"F7DE", x"F9C2", x"FA8A", x"F9BE", x"F94E", x"F944", x"F8A0", x"F8CF", x"FA0A", x"FA79", x"FAEC", x"FD26", x"FF2E", x"FFA3", x"FF87", x"FE5C", x"FB88", x"F9FE", x"FB64", x"FD4A", x"FF08", x"010F", x"0229", x"0233", x"0370", x"05AF", x"0720", x"083A", x"0914", x"088F", x"073E", x"0642", x"04EE", x"0365", x"02BA", x"0279", x"0224", x"025A", x"02D0", x"02C2", x"032A", x"045B", x"058E", x"06E0", x"0825", x"0817", x"06BF", x"04F9", x"0295", x"FFC8", x"FDE6", x"FC4A", x"FA64", x"F8EE", x"F7AF", x"F5B8", x"F485", x"F50D", x"F5A0", x"F588", x"F536", x"F36E", x"F068", x"EF3F", x"F0A8", x"F308", x"F66F", x"FA83", x"FD32", x"FEA0", x"0047", x"015B", x"016E", x"01BE", x"01C3", x"009F", x"FF18", x"FD76", x"FAC6", x"F7EC", x"F57F", x"F26D", x"EF22", x"ECF5", x"EB5D", x"EA61", x"EB5E", x"EDCC", x"F052", x"F378", x"F672", x"F7BA", x"F7B0", x"F746", x"F5D2", x"F448", x"F3CD", x"F38C", x"F359", x"F421", x"F50F", x"F565", x"F6E7", x"F8FC", x"F99E", x"F8D9", x"F726", x"F363", x"EFB7", x"EF3A", x"F0BB", x"F23E", x"F3F5", x"F4CD", x"F3B4", x"F2FC", x"F409", x"F544", x"F670", x"F7F3", x"F85E", x"F784", x"F6E4", x"F61D", x"F4FA", x"F495", x"F482", x"F3BA", x"F36F", x"F3F1", x"F45C", x"F582", x"F7CB", x"F976", x"FA7E", x"FBAF", x"FBB3", x"F9FC", x"F7E3", x"F4C9", x"F04D", x"EC88", x"EA18", x"E7E1", x"E702", x"E7D2", x"E81B", x"E86A", x"EA61", x"EC53", x"ED0B", x"EDCB", x"EDBF", x"EBE6", x"EB75", x"EDF8", x"F134", x"F48C", x"F82F", x"F9EF", x"F9AA", x"FA2D", x"FB71", x"FC5E", x"FDBB", x"FEE4", x"FDC1", x"FAED", x"F74F", x"F29D", x"EDED", x"EAD0", x"E823", x"E582", x"E3DE", x"E296", x"E13F", x"E15F", x"E2A9", x"E3F5", x"E633", x"E97D", x"EC33", x"EE40", x"F01A", x"F053", x"EF48", x"EF4B", x"F02D", x"F164", x"F3F0", x"F6D2", x"F843", x"F979", x"FBAB", x"FD46", x"FDCD", x"FDF1", x"FC5F", x"F904", x"F69E", x"F5FE", x"F5BD", x"F60B", x"F6F1", x"F73B", x"F731", x"F829", x"F9C3", x"FB34", x"FCC8", x"FDCA", x"FD6A", x"FBD9", x"F9AB", x"F710", x"F51D", x"F427", x"F3B2", x"F385", x"F38A", x"F346", x"F2D7", x"F2EA", x"F36E", x"F43A", x"F593", x"F6ED", x"F778", x"F75D", x"F6B2", x"F537", x"F397", x"F254", x"F12D", x"F05A", x"F080", x"F109", x"F164", x"F243", x"F34C", x"F336", x"F201", x"F026", x"ED8F", x"EB2C", x"EB32", x"ED9F", x"F11F", x"F513", x"F922", x"FC15", x"FDE1", x"FF54", x"0083", x"0115", x"016D", x"015E", x"FFFE", x"FCEA", x"F87E", x"F360", x"EE89", x"EA77", x"E75C", x"E56B", x"E4A9", x"E49C", x"E555", x"E6DD", x"E86A", x"EA06", x"EC37", x"EE89", x"F01C", x"F127", x"F178", x"F083", x"EF81", x"EF6E", x"EFDF", x"F118", x"F396", x"F619", x"F7F5", x"FA4F", x"FC83", x"FCC4", x"FBA2", x"F990", x"F5DE", x"F25D", x"F1AF", x"F26D", x"F2AA", x"F2EC", x"F2A7", x"F109", x"F02E", x"F18F", x"F38E", x"F5B6", x"F876", x"FA78", x"FABF", x"FA84", x"F9BB", x"F824", x"F711", x"F6BD", x"F649", x"F645", x"F6FA", x"F756", x"F7A0", x"F8C4", x"F9B0", x"FA78", x"FBE3", x"FCB3", x"FB89", x"F948", x"F630", x"F212", x"EEE1", x"ED90", x"ECF8", x"ED18", x"EE69", x"EF93", x"F092", x"F2D2", x"F537", x"F65B", x"F6DD", x"F6CD", x"F58A", x"F56D", x"F7F7", x"FB74", x"FF0E", x"02B2", x"04F8", x"055A", x"05AB", x"063A", x"0692", x"0777", x"08CB", x"093E", x"08D9", x"07B5", x"055C", x"0297", x"001D", x"FD2D", x"FA31", x"F829", x"F6A9", x"F5CA", x"F6AA", x"F822", x"F90E", x"FA55", x"FBE5", x"FC7E", x"FD05", x"FE21", x"FE1E", x"FD9B", x"FE5F", x"FF7A", x"005E", x"027C", x"04B2", x"0545", x"0620", x"0838", x"0951", x"095D", x"0944", x"0753", x"03C7", x"0202", x"021E", x"01FF", x"0232", x"02DB", x"0263", x"01CE", x"02F2", x"04BB", x"0641", x"085F", x"0A69", x"0B4B", x"0B95", x"0B65", x"09F4", x"080B", x"0676", x"049F", x"032A", x"02DE", x"031E", x"03D3", x"057C", x"0752", x"086C", x"0944", x"096B", x"081B", x"062F", x"044F", x"01F3", x"FFCA", x"FE76", x"FD22", x"FBD0", x"FB7F", x"FB98", x"FBA7", x"FCE9", x"FF24", x"003F", x"0054", x"FFD7", x"FE49", x"FCDF", x"FE5B", x"01E5", x"057F", x"0900", x"0C29", x"0DB3", x"0E63", x"0F89", x"1080", x"1107", x"120B", x"133B", x"134F", x"11EA", x"0EF6", x"0A8D", x"05C3", x"0160", x"FD6D", x"FA8F", x"F8C5", x"F7B2", x"F7C2", x"F936", x"FACA", x"FC98", x"FF45", x"0199", x"027D", x"0285", x"0160", x"FE92", x"FC50", x"FC13", x"FC88", x"FDD5", x"003E", x"01F6", x"02EA", x"0531", x"0815", x"0943", x"0946", x"07C8", x"03AA", x"FFA9", x"FEC8", x"FF79", x"0089", x"02B3", x"045F", x"046C", x"04F5", x"0691", x"0785", x"089F", x"0AC9", x"0C66", x"0D5A", x"0E6A", x"0E86", x"0D9E", x"0D55", x"0D48", x"0CDD", x"0D3F", x"0DF3", x"0DDB", x"0E4C", x"0FC8", x"1104", x"12DA", x"15F5", x"17C0", x"1761", x"15CE", x"123A", x"0CFF", x"091D", x"0725", x"05B7", x"05CF", x"0724", x"0799", x"0850", x"0ABD", x"0CFE", x"0E36", x"0F50", x"0E84", x"0BAC", x"0A65", x"0BC0", x"0E3F", x"12A3", x"1836", x"1C0F", x"1EA2", x"21D7", x"244F", x"257D", x"26AF", x"2688", x"23BA", x"205D", x"1CE8", x"1873", x"147F", x"11BF", x"0E92", x"0B77", x"09A4", x"07E0", x"05E5", x"0551", x"0567", x"05B4", x"074A", x"098A", x"0AA3", x"0B21", x"0B2A", x"09E1", x"08C5", x"0903", x"098F", x"0A91", x"0CBF", x"0E4E", x"0ED2", x"1076", x"12E7", x"14AD", x"164A", x"16BF", x"13B2", x"0EBE", x"0B16", x"0890", x"0751", x"0843", x"09D7", x"0A57", x"0AE9", x"0C27", x"0D0E", x"0E14", x"0FD5", x"115E", x"1231", x"1258", x"112B", x"0EA4", x"0BB3", x"08F8", x"0719", x"0695", x"0710", x"085A", x"0AB9", x"0D80", x"1035", x"12F2", x"14D5", x"14D1", x"1406", x"12DF", x"10D2", x"0E92", x"0D7C", x"0C86", x"0BDB", x"0CFF", x"0EC7", x"0EDC", x"0E40", x"0E29", x"0D8E", x"0CD9", x"0CF9", x"0BDB", x"080F", x"046C", x"033E", x"03C3", x"05E1", x"0992", x"0C99", x"0DAA", x"0E7F", x"0FE8", x"10F4", x"1200", x"1401", x"15D8", x"1678", x"15EB", x"13C2", x"0F8A", x"0A76", x"05C5", x"01C1", x"FEDA", x"FD8A", x"FD62", x"FE4E", x"004D", x"02AA", x"04C3", x"06BC", x"07BE", x"0733", x"05FF", x"04BF", x"039B", x"03D5", x"05BB", x"07E0", x"09A6", x"0B89", x"0CB6", x"0D7E", x"0F79", x"11AD", x"11C5", x"0FF5", x"0C79", x"06FC", x"0219", x"00C6", x"0155", x"022C", x"03FF", x"05D0", x"05E8", x"05F5", x"06F1", x"0714", x"06F6", x"089A", x"0B00", x"0C83", x"0D7A", x"0D72", x"0BAB", x"0962", x"07BA", x"0637", x"04CA", x"03C0", x"033E", x"0383", x"0490", x"05C1", x"0701", x"0810", x"081F", x"0771", x"067A", x"04B7", x"02B4", x"01C1", x"0193", x"01BA", x"02FB", x"0488", x"0560", x"06AF", x"08C0", x"0A01", x"0A77", x"0A31", x"078B", x"0367", x"010F", x"00E9", x"0239", x"05E5", x"0A5D", x"0D04", x"0EDE", x"1122", x"122B", x"11F7", x"11C5", x"103F", x"0D0F", x"0A95", x"0884", x"05A2", x"02F8", x"00B9", x"FD58", x"FA49", x"F902", x"F823", x"F781", x"F857", x"F97B", x"FA3A", x"FC24", x"FEBB", x"0026", x"0116", x"020E", x"023E", x"02BA", x"04CC", x"0741", x"0997", x"0C63", x"0EB2", x"103F", x"12CD", x"164C", x"196A", x"1C18", x"1D6A", x"1B6E", x"1766", x"13D8", x"10EC", x"0EE5", x"0ED7", x"0FB3", x"0FDE", x"1053", x"1173", x"11E2", x"11D0", x"126A", x"134B", x"1415", x"1561", x"1688", x"1641", x"14D0", x"132F", x"117C", x"1014", x"0F9E", x"1024", x"1137", x"130E", x"15C0", x"187F", x"1A31", x"1AAF", x"1A35", x"18C9", x"16ED", x"1596", x"1498", x"1349", x"1221", x"11C6", x"112D", x"0FD3", x"0EEB", x"0ECE", x"0F05", x"0FEC", x"1147", x"10B1", x"0D70", x"09EC", x"07D9", x"073C", x"08D2", x"0C78", x"0FD6", x"11EB", x"13E9", x"159D", x"15FC", x"160E", x"16BF", x"1747", x"1771", x"1792", x"1645", x"129E", x"0DF2", x"091F", x"047E", x"0144", x"FFE1", x"FF5C", x"FF90", x"0099", x"0184", x"01D7", x"01C9", x"00C7", x"FE94", x"FC4F", x"FA7C", x"F948", x"F97B", x"FAF3", x"FCC8", x"FF2D", x"01F6", x"042E", x"0697", x"09FE", x"0CEB", x"0E84", x"0F34", x"0D89", x"0959", x"05C3", x"0428", x"0312", x"02F0", x"041C", x"046C", x"03B5", x"040E", x"04A1", x"0401", x"03D6", x"047F", x"04C0", x"0504", x"0594", x"048C", x"01DA", x"FEEF", x"FBDA", x"F921", x"F86C", x"F93E", x"FA88", x"FCCD", x"FF51", x"00F6", x"0263", x"03D5", x"03EB", x"02E6", x"0175", x"FF2F", x"FCD8", x"FBF3", x"FBFE", x"FC7B", x"FDDC", x"FED1", x"FEA3", x"FECF", x"FFAC", x"003B", x"0153", x"027F", x"0168", x"FED2", x"FD49", x"FC83", x"FC7A", x"FED2", x"0220", x"043A", x"0659", x"08FD", x"0A3E", x"0A7C", x"0B24", x"0B29", x"0AA4", x"0AD0", x"0A8E", x"080E", x"042F", x"FF58", x"F9AA", x"F523", x"F303", x"F225", x"F21A", x"F2F6", x"F3AB", x"F3E4", x"F480", x"F50D", x"F4F9", x"F4E1", x"F4E3", x"F51C", x"F673", x"F8D3", x"FBC2", x"FF38", x"026D", x"03D6", x"0426", x"0489", x"04EE", x"0619", x"08D9", x"0AB7", x"09D9", x"07B2", x"0583", x"0334", x"0293", x"0418", x"0547", x"04FA", x"0477", x"0373", x"0165", x"FFC3", x"FF32", x"FEA1", x"FE64", x"FF04", x"FED2", x"FCFD", x"FA41", x"F6F1", x"F379", x"F16B", x"F139", x"F1F9", x"F364", x"F564", x"F748", x"F8A5", x"F98F", x"F99C", x"F893", x"F6F4", x"F54C", x"F408", x"F378", x"F358", x"F380", x"F3C4", x"F358", x"F1C7", x"F025", x"EF5D", x"EF83", x"F0FB", x"F342", x"F3EB", x"F1DA", x"EF00", x"ECC7", x"EBCE", x"ED77", x"F1D9", x"F677", x"FA14", x"FD57", x"FF75", x"FFBE", x"FFAA", x"FFFC", x"FFEB", x"FF8D", x"FF11", x"FCD2", x"F834", x"F276", x"EC73", x"E6BA", x"E2C0", x"E0CB", x"DFDB", x"DFB6", x"E06F", x"E157", x"E20E", x"E292", x"E272", x"E157", x"DFD8", x"DE6F", x"DDAE", x"DDD8", x"DF02", x"E153", x"E4A7", x"E7F0", x"EAC1", x"ED96", x"F01F", x"F1FB", x"F3E6", x"F50C", x"F382", x"EFE5", x"EC64", x"E946", x"E774", x"E846", x"EA5A", x"EB51", x"EBE7", x"EC73", x"EBE7", x"EB0C", x"EB42", x"EBA1", x"EBFD", x"EDAF", x"EFB9", x"F080", x"F075", x"EF96", x"ED44", x"EB1E", x"EAA0", x"EB19", x"EC3C", x"EE93", x"F0FB", x"F293", x"F3CA", x"F40E", x"F282", x"EFE7", x"ED3F", x"EACD", x"E9A3", x"E9E6", x"EADD", x"EC30", x"ED8D", x"EDDE", x"ED6A", x"ED2B", x"ED1D", x"ED79", x"EEFC", x"F01C", x"EF27", x"ECFD", x"EADB", x"E924", x"E96E", x"ECA2", x"F0D6", x"F48B", x"F80F", x"FAC6", x"FC1D", x"FCF6", x"FDC6", x"FDDC", x"FD81", x"FD3E", x"FC4B", x"FA13", x"F6D1", x"F2AC", x"EDF2", x"E9AB", x"E6A2", x"E4DD", x"E43B", x"E48C", x"E59F", x"E6C9", x"E738", x"E702", x"E657", x"E56C", x"E4E1", x"E5E1", x"E7F4", x"EA3D", x"ED3E", x"F0CC", x"F384", x"F552", x"F70B", x"F83D", x"F8F4", x"FA7B", x"FC5D", x"FC85", x"FAD1", x"F856", x"F571", x"F363", x"F3DA", x"F633", x"F887", x"FA43", x"FB42", x"FB0C", x"FA0A", x"F968", x"F925", x"F917", x"F9B2", x"FAED", x"FBD9", x"FBF7", x"FB66", x"FA31", x"F88E", x"F76B", x"F764", x"F7CA", x"F887", x"F9F3", x"FBA3", x"FCA4", x"FCED", x"FC30", x"F9F6", x"F70A", x"F504", x"F432", x"F425", x"F4C4", x"F582", x"F584", x"F4D4", x"F428", x"F3C5", x"F3C6", x"F489", x"F5D7", x"F711", x"F753", x"F692", x"F54F", x"F454", x"F43C", x"F5C5", x"F8C5", x"FC05", x"FEFE", x"01B4", x"03BB", x"04D8", x"05D2", x"06AA", x"06E2", x"06EB", x"06E7", x"0597", x"029A", x"FE8E", x"F980", x"F41B", x"F021", x"EDFD", x"ECDE", x"ECDC", x"EE0A", x"EF59", x"F050", x"F102", x"F0CD", x"EF36", x"ED64", x"EC51", x"EC54", x"ED6C", x"EFA3", x"F266", x"F4DE", x"F69D", x"F7DE", x"F8F3", x"F9CE", x"FAFB", x"FD04", x"FE82", x"FE2B", x"FC59", x"F9C1", x"F695", x"F4C0", x"F599", x"F77E", x"F939", x"FB3C", x"FCCC", x"FCDD", x"FCC0", x"FCF1", x"FC53", x"FBBF", x"FCCD", x"FE78", x"FF74", x"003F", x"0015", x"FE4D", x"FCC9", x"FCB9", x"FD4B", x"FE14", x"FF66", x"0078", x"00D4", x"00DF", x"0055", x"FEA5", x"FC38", x"F9D3", x"F7F7", x"F720", x"F717", x"F7D3", x"F93D", x"FA9C", x"FB77", x"FC35", x"FCFF", x"FD8D", x"FEEF", x"010A", x"0234", x"0180", x"FFD1", x"FD47", x"FB0E", x"FB53", x"FE54", x"0235", x"064C", x"09F7", x"0BE1", x"0C38", x"0C16", x"0B81", x"0A5A", x"0983", x"0905", x"0811", x"0670", x"040C", x"00B0", x"FD06", x"F9AE", x"F72C", x"F596", x"F4E9", x"F4E4", x"F5DF", x"F741", x"F7EE", x"F7CE", x"F728", x"F588", x"F3BA", x"F303", x"F2FB", x"F346", x"F515", x"F853", x"FB6A", x"FE25", x"00C9", x"0211", x"0263", x"036B", x"0487", x"0434", x"02CE", x"00AA", x"FD82", x"FB0C", x"FB18", x"FCD8", x"FF1C", x"0195", x"031A", x"028A", x"00DF", x"FF28", x"FD74", x"FC53", x"FCB9", x"FDEC", x"FEF7", x"FF69", x"FF02", x"FD33", x"FAD0", x"F935", x"F88A", x"F8B6", x"F9BC", x"FB5A", x"FCF2", x"FE46", x"FF44", x"FF52", x"FDDD", x"FB7E", x"F8EF", x"F6C5", x"F592", x"F5BE", x"F6D8", x"F813", x"F92B", x"F9C8", x"F9C6", x"F964", x"F933", x"F960", x"F99C", x"F969", x"F87D", x"F6DB", x"F4EC", x"F3D9", x"F47E", x"F6B2", x"F9BF", x"FD26", x"FFE6", x"0148", x"018A", x"012C", x"003B", x"FF34", x"FEEE", x"FEF5", x"FE8D", x"FD88", x"FBBC", x"F8EA", x"F5ED", x"F3BF", x"F242", x"F15B", x"F13A", x"F1B7", x"F2A2", x"F3EF", x"F567", x"F657", x"F66E", x"F5B4", x"F4B3", x"F3DD", x"F36A", x"F3C9", x"F54D", x"F739", x"F920", x"FB14", x"FC81", x"FCE9", x"FDAD", x"FF54", x"005C", x"0039", x"FF44", x"FC7B", x"F8DB", x"F7AA", x"F993", x"FC99", x"008D", x"049D", x"062D", x"057F", x"04B0", x"0318", x"0070", x"FF27", x"FFA1", x"0042", x"013E", x"0281", x"01F7", x"000D", x"FEC8", x"FE29", x"FDDB", x"FED5", x"0053", x"014E", x"0244", x"035D", x"0396", x"034D", x"02B8", x"013D", x"FF77", x"FE52", x"FDDB", x"FE58", x"0059", x"028E", x"0438", x"057E", x"0616", x"061C", x"072C", x"0921", x"0A6A", x"0AE9", x"0A26", x"074A", x"041C", x"0327", x"0427", x"065F", x"0A0F", x"0D6E", x"0EEB", x"0F8B", x"0FE9", x"0F00", x"0D6B", x"0C21", x"0A7B", x"084E", x"063B", x"03E9", x"013B", x"FEEF", x"FD03", x"FB26", x"F997", x"F836", x"F745", x"F7D3", x"F994", x"FB8D", x"FDEE", x"005A", x"01C5", x"02FB", x"04A4", x"05C8", x"0690", x"0896", x"0AF9", x"0CF9", x"0F90", x"121B", x"1322", x"141A", x"160F", x"1769", x"17ED", x"186B", x"1761", x"1491", x"1328", x"142F", x"1647", x"19AF", x"1DC0", x"1FA8", x"1F27", x"1E42", x"1CDE", x"1A8B", x"18B5", x"17DE", x"171B", x"16E9", x"17BE", x"1878", x"1892", x"18AD", x"18DD", x"1907", x"196E", x"1A41", x"1B70", x"1D11", x"1EC9", x"2004", x"2044", x"1F0C", x"1CA3", x"1A13", x"1831", x"170F", x"174C", x"18BE", x"1A48", x"1B6D", x"1C41", x"1C3A", x"1B64", x"1B0D", x"1B63", x"1B61", x"1AAA", x"1907", x"15C8", x"11E4", x"0FE7", x"10A9", x"139F", x"1863", x"1DD0", x"2201", x"2470", x"25FC", x"2689", x"25E8", x"24FA", x"2452", x"237C", x"2270", x"2137", x"1F9E", x"1D59", x"1AF2", x"18B1", x"1672", x"1406", x"119A", x"0FE3", x"0EE9", x"0E5B", x"0E1C", x"0DFA", x"0D2A", x"0C15", x"0B97", x"0B77", x"0B2C", x"0B93", x"0CDC", x"0E24", x"0FDA", x"1267", x"1469", x"15BB", x"1801", x"1AA6", x"1C53", x"1D40", x"1D24", x"1A9E", x"179F", x"16E7", x"17E6", x"19F0", x"1D51", x"203E", x"20E0", x"2078", x"1FB2", x"1D85", x"1ABA", x"189A", x"167E", x"1488", x"13F3", x"13DD", x"1357", x"130D", x"1272", x"10C9", x"0F3B", x"0E5A", x"0D66", x"0CED", x"0D41", x"0CC6", x"0B7E", x"0A87", x"095C", x"07F0", x"0780", x"07E5", x"0843", x"09A1", x"0BFB", x"0DF9", x"0FDB", x"11C5", x"12AF", x"1332", x"14A6", x"1615", x"16BE", x"1718", x"15E0", x"12B6", x"101F", x"0FB3", x"10DF", x"1439", x"1936", x"1D26", x"1F3E", x"2082", x"2075", x"1F0B", x"1DFD", x"1D4F", x"1C3F", x"1BA6", x"1B6F", x"1A87", x"1927", x"17B5", x"151B", x"11D0", x"0EE8", x"0C6E", x"0AA4", x"0AA4", x"0B8B", x"0C64", x"0D79", x"0E42", x"0E37", x"0E43", x"0EDA", x"0F62", x"1093", x"1294", x"141D", x"1569", x"173B", x"185A", x"1895", x"19AC", x"1B3D", x"1C56", x"1E21", x"200E", x"1F7A", x"1D32", x"1BBF", x"1AFE", x"1B23", x"1D8E", x"206A", x"212B", x"20B5", x"1FF8", x"1DF8", x"1B08", x"187F", x"15BE", x"12DB", x"1169", x"1188", x"123E", x"1378", x"14DB", x"1568", x"153D", x"14B3", x"13BC", x"12AD", x"11FD", x"1175", x"111C", x"10EE", x"103B", x"0ED8", x"0D12", x"0AC1", x"0822", x"0646", x"053E", x"046D", x"046E", x"0526", x"0524", x"04AA", x"04F6", x"058A", x"05F0", x"06E1", x"0759", x"0579", x"0297", x"0149", x"01AA", x"03DD", x"0873", x"0DA3", x"1107", x"12FA", x"1425", x"1366", x"110E", x"0E96", x"0C67", x"0A47", x"08DD", x"07E4", x"063A", x"03DE", x"012C", x"FE49", x"FB4B", x"F871", x"F5D5", x"F3FD", x"F2C4", x"F1AD", x"F0D0", x"F033", x"EF5E", x"EEC7", x"EF3C", x"EFC7", x"F03D", x"F1A7", x"F3E4", x"F61F", x"F91C", x"FC86", x"FE6A", x"FF8F", x"01BF", x"0443", x"06A2", x"099A", x"0B2C", x"096C", x"069B", x"04EE", x"03EE", x"046F", x"0715", x"0937", x"0986", x"0981", x"08FB", x"06F8", x"04D0", x"02F8", x"008D", x"FE9C", x"FE00", x"FDC4", x"FDE4", x"FED4", x"FF17", x"FE80", x"FE27", x"FDCB", x"FD20", x"FDB3", x"FEBA", x"FE8B", x"FE13", x"FDEC", x"FCC0", x"FB36", x"FA5E", x"F8F2", x"F6EA", x"F64E", x"F6AA", x"F700", x"F833", x"F9B5", x"FA0C", x"FA8B", x"FBFF", x"FD0B", x"FD8C", x"FDEF", x"FC62", x"F90E", x"F6BE", x"F63C", x"F77A", x"FB97", x"0129", x"0558", x"07C0", x"0912", x"0860", x"06C2", x"05B5", x"047A", x"02B1", x"0174", x"FFFC", x"FDBF", x"FBCF", x"FA01", x"F739", x"F489", x"F28D", x"F050", x"EE82", x"EE00", x"ED78", x"ECBE", x"ED01", x"EDA2", x"EDF5", x"EED1", x"EFF4", x"F06F", x"F179", x"F387", x"F57F", x"F7C8", x"FA6D", x"FBB6", x"FBA2", x"FBEF", x"FC45", x"FCCA", x"FEF7", x"017A", x"0192", x"004B", x"FF0C", x"FD88", x"FD5B", x"FFFE", x"031D", x"049D", x"0591", x"05C3", x"0429", x"023B", x"00B7", x"FE66", x"FBF9", x"FAFA", x"FADF", x"FAEC", x"FBCA", x"FC9D", x"FC7A", x"FC4D", x"FC91", x"FC97", x"FCC5", x"FD4B", x"FD47", x"FCAC", x"FBE4", x"FA4F", x"F7D8", x"F526", x"F246", x"EF6E", x"EDE2", x"ED9D", x"EE39", x"F02B", x"F2D2", x"F45C", x"F50F", x"F58F", x"F567", x"F50D", x"F5B5", x"F5D1", x"F40B", x"F210", x"F170", x"F200", x"F4F6", x"FA6D", x"FFA2", x"02F5", x"055C", x"0673", x"05DE", x"04D8", x"03FE", x"029C", x"015D", x"00F7", x"0087", x"FFD6", x"FF17", x"FD6A", x"FA8D", x"F726", x"F33B", x"EF5F", x"ECF9", x"EC0A", x"EBD0", x"EC71", x"ED5C", x"ED4F", x"ED11", x"ED4D", x"ED10", x"ECDA", x"EDCF", x"EEEF", x"EFC2", x"F16D", x"F2D4", x"F28A", x"F22A", x"F2ED", x"F39B", x"F51E", x"F7B9", x"F8C0", x"F73C", x"F5EF", x"F585", x"F61B", x"F93C", x"FE21", x"0180", x"02DF", x"032F", x"0182", x"FEA5", x"FC99", x"FB09", x"F991", x"F961", x"FA05", x"FA79", x"FB88", x"FCFA", x"FD46", x"FCBA", x"FBF9", x"FA24", x"F817", x"F72A", x"F645", x"F4B5", x"F345", x"F166", x"EE72", x"EBDC", x"E9E8", x"E7C1", x"E656", x"E62A", x"E5FE", x"E63D", x"E78A", x"E8A8", x"E94D", x"EADE", x"EC90", x"EDAC", x"EF67", x"F0FE", x"F09C", x"EF43", x"EE7F", x"EE13", x"EF55", x"F37E", x"F8A9", x"FCE3", x"0086", x"02A7", x"0291", x"01E7", x"0140", x"FFBC", x"FE53", x"FDAF", x"FCDE", x"FBFB", x"FBED", x"FB3E", x"F938", x"F6E4", x"F421", x"F097", x"EDB1", x"EBF2", x"EA59", x"E97E", x"E9E9", x"EA9C", x"EB71", x"ECAC", x"ED8B", x"EDC7", x"EE63", x"EEF7", x"EF21", x"EFFF", x"F13E", x"F1DD", x"F2A5", x"F406", x"F4EB", x"F5F8", x"F82E", x"F9C6", x"F954", x"F80F", x"F65F", x"F46F", x"F440", x"F69F", x"F972", x"FB9F", x"FD4F", x"FD94", x"FC0E", x"F9EB", x"F7A9", x"F51B", x"F355", x"F2FE", x"F370", x"F45C", x"F581", x"F5CF", x"F529", x"F3E5", x"F244", x"F074", x"EF41", x"EEC8", x"EEA7", x"EEEA", x"EED7", x"EDCA", x"EBE4", x"E98C", x"E730", x"E5E4", x"E610", x"E6F6", x"E85C", x"EA67", x"EBD8", x"EC34", x"EC57", x"EC39", x"EB61", x"EB2E", x"EBEE", x"EB99", x"E9B7", x"E7C1", x"E5F2", x"E4DA", x"E64F", x"E9FC", x"ED3B", x"EF99", x"F179", x"F210", x"F183", x"F119", x"F0AB", x"EFA7", x"EF1B", x"EF26", x"EF32", x"EF65", x"EFC2", x"EF4F", x"EE17", x"EC6E", x"E9FC", x"E729", x"E51D", x"E3BF", x"E2EA", x"E33A", x"E425", x"E4BA", x"E542", x"E5A0", x"E525", x"E485", x"E46B", x"E47B", x"E50C", x"E6BD", x"E87B", x"E9CF", x"EB9B", x"EDA3", x"EF7D", x"F23A", x"F547", x"F67A", x"F5CC", x"F471", x"F272", x"F11A", x"F290", x"F5D3", x"F8F9", x"FBC6", x"FD9B", x"FD24", x"FB44", x"F94C", x"F71A", x"F553", x"F502", x"F58B", x"F640", x"F745", x"F7F2", x"F7CB", x"F770", x"F6F3", x"F5F3", x"F508", x"F45C", x"F363", x"F2B1", x"F297", x"F26D", x"F20D", x"F1CC", x"F0DB", x"EF5E", x"EE56", x"EDC1", x"ED7B", x"EEA5", x"F0C1", x"F2A5", x"F4A1", x"F6A3", x"F78F", x"F81F", x"F9A6", x"FAC0", x"FA8E", x"F9F1", x"F891", x"F663", x"F5DA", x"F7FB", x"FAFB", x"FE05", x"00EB", x"01F1", x"00FA", x"FFAF", x"FE4F", x"FC5D", x"FAC2", x"F9F2", x"F92D", x"F891", x"F879", x"F827", x"F76D", x"F6B7", x"F5D5", x"F46E", x"F2AC", x"F0A8", x"EEF5", x"EE45", x"EEB0", x"EFD3", x"F196", x"F30F", x"F41D", x"F587", x"F73C", x"F883", x"F9B8", x"FB16", x"FBBE", x"FBEE", x"FCC5", x"FDCA", x"FEC8", x"0114", x"045B", x"06C4", x"079E", x"0736", x"0517", x"0276", x"01C2", x"0324", x"0523", x"070D", x"083B", x"078A", x"0528", x"0257", x"FF5A", x"FC2D", x"F9D6", x"F8F3", x"F90B", x"F995", x"FA9D", x"FBD2", x"FCC2", x"FDC8", x"FF13", x"FFF3", x"FFC3", x"FF75", x"FFAF", x"003B", x"00CE", x"0146", x"00A2", x"FE85", x"FC60", x"FB7E", x"FB71", x"FC13", x"FDBB", x"FFA0", x"00A8", x"012D", x"017D", x"0107", x"004A", x"00B2", x"01EA", x"023D", x"0159", x"FFAA", x"FD51", x"FB87", x"FC63", x"FFAE", x"03A8", x"0773", x"0AD0", x"0C5A", x"0C00", x"0AFA", x"09AD", x"0819", x"075F", x"0802", x"08A7", x"0876", x"0793", x"05DA", x"0345", x"0100", x"FF71", x"FDA1", x"FB73", x"F97D", x"F7FD", x"F6DB", x"F662", x"F692", x"F696", x"F640", x"F633", x"F6BB", x"F709", x"F72C", x"F7CA", x"F872", x"F865", x"F861", x"F8BF", x"F8EF", x"F9BB", x"FCBB", x"00BE", x"0395", x"056F", x"0650", x"05C2", x"0556", x"070D", x"09B5", x"0BA9", x"0D53", x"0E2F", x"0D04", x"0ABA", x"088C", x"05F4", x"034D", x"01DA", x"010F", x"0011", x"FEEE", x"FDD5", x"FC7F", x"FB92", x"FB75", x"FB91", x"FB2D", x"FA53", x"F906", x"F7DA", x"F733", x"F71D", x"F738", x"F701", x"F619", x"F4FC", x"F41B", x"F348", x"F2F0", x"F3A1", x"F49D", x"F563", x"F689", x"F7B6", x"F875", x"F9DF", x"FCCE", x"FF8C", x"0117", x"01D1", x"0168", x"0033", x"00A3", x"03A9", x"078F", x"0B45", x"0E92", x"107B", x"10AB", x"106A", x"103F", x"0FB6", x"0EFC", x"0E93", x"0E0F", x"0CC2", x"0AD6", x"08C7", x"06BA", x"04AE", x"02F3", x"0165", x"FF5D", x"FD28", x"FC09", x"FC18", x"FCA2", x"FDA7", x"FEC0", x"FEDD", x"FEA7", x"FF67", x"009C", x"01AC", x"0369", x"056E", x"069C", x"07AB", x"093C", x"0A12", x"0A81", x"0C54", x"0F0C", x"1124", x"12BA", x"1365", x"120E", x"1001", x"0FCC", x"111C", x"12A6", x"1441", x"1553", x"14BC", x"12F5", x"1176", x"1020", x"0EA6", x"0DE4", x"0E43", x"0EB1", x"0E47", x"0D64", x"0C2F", x"0AAF", x"09AB", x"09AB", x"0994", x"0897", x"0786", x"0718", x"06ED", x"06E2", x"0705", x"064D", x"0461", x"0275", x"014A", x"008C", x"0096", x"01D6", x"0392", x"050F", x"063E", x"06E4", x"064A", x"054D", x"0513", x"057E", x"05D2", x"05F9", x"05D4", x"0529", x"0509", x"0707", x"0ACC", x"0EC1", x"1278", x"153C", x"15B0", x"13F7", x"11AD", x"0F48", x"0CD8", x"0BE9", x"0CC9", x"0D25", x"0BBF", x"0922", x"053E", x"005D", x"FC3D", x"F995", x"F6B8", x"F397", x"F187", x"F0C9", x"F0CE", x"F1F2", x"F3D5", x"F528", x"F5B3", x"F69F", x"F7DE", x"F8C6", x"F9C0", x"FB5D", x"FD0C", x"FE5F", x"0017", x"0234", x"043E", x"06FB", x"0AFF", x"0EC7", x"10B4", x"1109", x"0FD3", x"0D6C", x"0BFD", x"0D14", x"0F67", x"11B1", x"13FB", x"152C", x"1483", x"1346", x"1250", x"10E4", x"0F5B", x"0ED3", x"0E7E", x"0D78", x"0C32", x"0AFD", x"098E", x"08D5", x"0953", x"0A2C", x"0A26", x"093D", x"07FE", x"06E1", x"0670", x"06EC", x"0829", x"0929", x"097E", x"09A5", x"0991", x"08D4", x"083E", x"08AF", x"0974", x"09E8", x"0AB4", x"0B4A", x"0B19", x"0B97", x"0D97", x"0F76", x"106F", x"111C", x"10EA", x"0FF2", x"105E", x"129C", x"1503", x"170A", x"18E6", x"1954", x"1826", x"16C9", x"1579", x"13C0", x"1296", x"1278", x"128D", x"1227", x"1181", x"1081", x"0F1D", x"0DE1", x"0D20", x"0C16", x"0A2A", x"07B5", x"0586", x"03E0", x"030A", x"0347", x"0434", x"04B3", x"04FE", x"0589", x"05AA", x"0550", x"05C6", x"072B", x"0896", x"0A8B", x"0CF0", x"0E8B", x"0FA8", x"120F", x"1560", x"1807", x"19E5", x"1A4B", x"183E", x"152C", x"1396", x"138D", x"144A", x"15D3", x"1734", x"171D", x"15D8", x"1477", x"1346", x"12A3", x"135F", x"1524", x"16D9", x"1772", x"16E1", x"1591", x"140D", x"12E1", x"1268", x"121E", x"114A", x"0FFC", x"0EE3", x"0DDD", x"0CBE", x"0BFC", x"0B33", x"09C5", x"083B", x"0740", x"068C", x"0674", x"07E7", x"0A33", x"0C4D", x"0E59", x"0FDB", x"1024", x"102C", x"1172", x"133B", x"1490", x"157E", x"152E", x"1326", x"1156", x"119A", x"1369", x"15E1", x"18FC", x"1B53", x"1BB6", x"1ACA", x"199B", x"17EB", x"165E", x"1601", x"16A0", x"16C9", x"1628", x"14B8", x"1263", x"0FA7", x"0D3C", x"0B2B", x"08DB", x"063E", x"040F", x"02AA", x"024D", x"02FD", x"0472", x"05D5", x"0694", x"06BA", x"0671", x"05B5", x"052C", x"050D", x"04F8", x"0500", x"0566", x"05F9", x"06AA", x"0850", x"0AC6", x"0CF4", x"0E8E", x"0F4D", x"0E41", x"0C2E", x"0B47", x"0C3D", x"0E2C", x"10E1", x"1374", x"142A", x"1316", x"11B7", x"1022", x"0E4F", x"0D28", x"0CFC", x"0CEB", x"0C8B", x"0C05", x"0AF8", x"09D5", x"0942", x"095F", x"09C5", x"09E1", x"096F", x"08B7", x"0850", x"081B", x"0823", x"08A2", x"08D1", x"07F2", x"0646", x"03A9", x"0007", x"FC7A", x"FA3B", x"F8C1", x"F807", x"F823", x"F83A", x"F817", x"F937", x"FBB1", x"FE56", x"0114", x"034C", x"036F", x"0271", x"02B6", x"044C", x"0688", x"09E6", x"0D76", x"0F38", x"0FC8", x"102D", x"0F72", x"0D70", x"0BDA", x"0B17", x"0A72", x"0A5B", x"0AF5", x"0B47", x"0B56", x"0BE2", x"0CBF", x"0D02", x"0C41", x"0ABA", x"08CD", x"06D3", x"053A", x"045C", x"03BF", x"02BA", x"0163", x"0005", x"FE2F", x"FC62", x"FBCE", x"FC4C", x"FD36", x"FEB8", x"003B", x"00BB", x"0123", x"02A6", x"04C4", x"0718", x"09C6", x"0B34", x"0A55", x"08BE", x"07BC", x"0714", x"0771", x"0908", x"09D9", x"0929", x"0813", x"06CB", x"0516", x"03F4", x"03B0", x"032C", x"0265", x"018E", x"003C", x"FE7E", x"FD23", x"FBEE", x"FAD6", x"F9FB", x"F90D", x"F7F0", x"F74C", x"F6CF", x"F5FC", x"F54E", x"F4CD", x"F3C1", x"F2D1", x"F286", x"F222", x"F1E4", x"F2C3", x"F3F6", x"F487", x"F4F9", x"F4DE", x"F397", x"F299", x"F30E", x"F3F5", x"F4CA", x"F59C", x"F4D4", x"F256", x"F05A", x"F022", x"F10F", x"F38B", x"F6D9", x"F8B2", x"F883", x"F79F", x"F5F4", x"F3B2", x"F244", x"F22B", x"F27C", x"F33F", x"F423", x"F3F1", x"F205", x"EF32", x"EBE1", x"E851", x"E520", x"E29F", x"E0BF", x"DFAC", x"DFA9", x"E0A6", x"E22D", x"E37B", x"E47C", x"E558", x"E5D0", x"E61A", x"E6C7", x"E796", x"E819", x"E933", x"EB1F", x"ECA6", x"EDEB", x"EFD8", x"F1A1", x"F2F6", x"F495", x"F5A7", x"F43D", x"F1B0", x"EFF1", x"EF20", x"EFD1", x"F2E7", x"F69F", x"F8EA", x"FA64", x"FB6B", x"FB10", x"F9EC", x"F916", x"F7E3", x"F642", x"F524", x"F443", x"F302", x"F211", x"F180", x"F0EF", x"F07C", x"F039", x"EF92", x"EEE2", x"EEA8", x"EECD", x"EF93", x"F14A", x"F314", x"F477", x"F598", x"F5A8", x"F471", x"F310", x"F1E4", x"F08B", x"EFEF", x"F02A", x"EFC1", x"EF2E", x"F030", x"F22F", x"F494", x"F7E0", x"FAA0", x"FAA5", x"F98A", x"F964", x"F9A3", x"FA65", x"FC95", x"FE96", x"FEC4", x"FE37", x"FD72", x"FB2F", x"F82A", x"F5E9", x"F42D", x"F2D5", x"F26C", x"F286", x"F25C", x"F24B", x"F295", x"F2E7", x"F339", x"F328", x"F2B6", x"F228", x"F181", x"F097", x"EFC8", x"EF11", x"EDF8", x"ECF1", x"EC75", x"EBFE", x"EBED", x"ED08", x"EEA9", x"F05F", x"F2C2", x"F50A", x"F65A", x"F807", x"FABD", x"FDCD", x"0186", x"05F1", x"0868", x"07FC", x"0651", x"03D2", x"00BF", x"FEE9", x"FE76", x"FD94", x"FC64", x"FBF4", x"FB3F", x"FA67", x"FA69", x"FA8E", x"FA2D", x"FA04", x"F9F0", x"F931", x"F8B4", x"F890", x"F7D4", x"F740", x"F7B2", x"F849", x"F941", x"FB55", x"FD04", x"FD52", x"FD58", x"FCED", x"FB42", x"F97E", x"F869", x"F744", x"F6F1", x"F859", x"FA50", x"FC41", x"FE58", x"FF7A", x"FF34", x"FF12", x"FF4A", x"FF9D", x"0125", x"0342", x"03C0", x"02E6", x"0233", x"0153", x"0106", x"02C8", x"04F0", x"0573", x"0500", x"0408", x"01A3", x"FF27", x"FDFA", x"FD83", x"FDBA", x"FF49", x"0112", x"0196", x"00E6", x"FEE3", x"FB8D", x"F815", x"F567", x"F372", x"F279", x"F28D", x"F2F1", x"F3A1", x"F49A", x"F542", x"F59F", x"F5ED", x"F5D9", x"F575", x"F550", x"F4E4", x"F431", x"F43E", x"F4E5", x"F543", x"F60B", x"F74E", x"F7DD", x"F867", x"F9D5", x"FA66", x"F909", x"F765", x"F651", x"F595", x"F718", x"FB0F", x"FEDA", x"0118", x"02BC", x"031C", x"019C", x"FFC0", x"FDFB", x"FB97", x"F934", x"F794", x"F5E2", x"F3C2", x"F1BD", x"EFBB", x"EDCC", x"EC87", x"EBFC", x"EBF5", x"ECE7", x"EE84", x"F044", x"F247", x"F434", x"F51A", x"F545", x"F4E2", x"F35B", x"F0FD", x"EF05", x"ED2B", x"EB64", x"EAA7", x"EA5C", x"E968", x"E8BC", x"E952", x"EA93", x"ECEE", x"F0CD", x"F3D1", x"F485", x"F449", x"F3CB", x"F2FF", x"F386", x"F5FB", x"F85E", x"FA2F", x"FC46", x"FD8F", x"FCF8", x"FBAE", x"F9E6", x"F74D", x"F524", x"F44A", x"F3E7", x"F3EE", x"F49C", x"F522", x"F54D", x"F5B8", x"F5EB", x"F5CA", x"F5FF", x"F603", x"F564", x"F517", x"F566", x"F5A0", x"F64E", x"F7A1", x"F861", x"F8ED", x"FA33", x"FB8D", x"FCA7", x"FE3E", x"FF80", x"FFC8", x"002D", x"011A", x"01C3", x"032B", x"0528", x"05C1", x"04F8", x"03FD", x"026D", x"0107", x"0180", x"02E5", x"0377", x"040D", x"048E", x"03C5", x"02D8", x"02BD", x"020B", x"00F9", x"0115", x"0143", x"00EE", x"012E", x"00F9", x"FEF0", x"FC8E", x"FAE9", x"F936", x"F892", x"F98D", x"FA2F", x"F9C0", x"F979", x"F8A2", x"F6F4", x"F5C9", x"F52F", x"F470", x"F4B6", x"F62F", x"F799", x"F94A", x"FB28", x"FBCC", x"FBAD", x"FBEA", x"FBC8", x"FBE5", x"FDC2", x"FF9D", x"FF70", x"FE57", x"FC74", x"F955", x"F7A3", x"F8C7", x"FA15", x"FAA3", x"FB82", x"FB58", x"F986", x"F85D", x"F7D7", x"F681", x"F5DC", x"F6DC", x"F7CE", x"F832", x"F84C", x"F65C", x"F1EB", x"ECF8", x"E83E", x"E3D9", x"E0F2", x"DF93", x"DEAC", x"DE6F", x"DEF6", x"DF85", x"E048", x"E165", x"E25F", x"E3A2", x"E58D", x"E749", x"E930", x"EC25", x"EF3F", x"F1F6", x"F525", x"F821", x"F9BD", x"FBC1", x"FE9B", x"0010", x"FFB1", x"FEDF", x"FD0E", x"FAE4", x"FB37", x"FDD8", x"0057", x"0273", x"0472", x"04BD", x"0385", x"023A", x"009E", x"FE53", x"FCBD", x"FC2D", x"FBB8", x"FB65", x"FB12", x"FA08", x"F877", x"F70B", x"F5BF", x"F4E1", x"F4DF", x"F534", x"F5B1", x"F667", x"F6F5", x"F71F", x"F773", x"F7B5", x"F76C", x"F70D", x"F6A2", x"F596", x"F4B7", x"F4DC", x"F538", x"F5C7", x"F76F", x"F9BB", x"FC42", x"0043", x"0559", x"08EB", x"0A8B", x"0AFB", x"09A3", x"0763", x"067A", x"06B6", x"0655", x"05F8", x"05E2", x"0473", x"01CE", x"FEFD", x"FB84", x"F7A3", x"F53A", x"F49E", x"F4E1", x"F632", x"F7C9", x"F82D", x"F79E", x"F6EA", x"F5E4", x"F544", x"F5E5", x"F6AB", x"F6C2", x"F6D3", x"F660", x"F4DD", x"F35D", x"F243", x"F0E2", x"F042", x"F10C", x"F249", x"F3D0", x"F5F7", x"F79F", x"F8D0", x"FABB", x"FD4E", x"005C", x"04F6", x"0A19", x"0D55", x"0EDB", x"0EF0", x"0CD7", x"0A4E", x"0963", x"08CB", x"07A2", x"074D", x"0710", x"05C4", x"04CD", x"0464", x"02D2", x"0116", x"00AA", x"0070", x"0056", x"0138", x"0195", x"007C", x"FF95", x"FF31", x"FEE4", x"FFF9", x"0250", x"03BF", x"044B", x"048B", x"0381", x"0186", x"FFFB", x"FE42", x"FC47", x"FB8A", x"FBB3", x"FC2E", x"FDDD", x"0038", x"01EB", x"03D4", x"05F9", x"0728", x"08A4", x"0BAA", x"0E02", x"0EE1", x"0F84", x"0EEF", x"0D2B", x"0DAD", x"1097", x"12FB", x"14B8", x"1626", x"1511", x"120D", x"0FD2", x"0D84", x"0A7F", x"0911", x"0963", x"09C6", x"0A82", x"0B17", x"094A", x"055D", x"013C", x"FD14", x"FA15", x"F9BA", x"FB33", x"FD25", x"FFCC", x"021F", x"0366", x"0480", x"05AC", x"05F7", x"0628", x"06AA", x"0669", x"062A", x"06C3", x"0707", x"06A7", x"06CC", x"0697", x"05C4", x"0668", x"0879", x"09CA", x"0A73", x"0AC6", x"0991", x"083B", x"0982", x"0CA8", x"0FDC", x"1389", x"16BE", x"17E2", x"177B", x"167B", x"13F7", x"105A", x"0D6C", x"0B53", x"09BA", x"08D7", x"07F4", x"0667", x"047F", x"02B2", x"011D", x"00B0", x"019F", x"0363", x"05BB", x"0824", x"092D", x"0909", x"087E", x"0769", x"05EE", x"04EE", x"03F3", x"022A", x"0089", x"FF46", x"FDA3", x"FC3F", x"FC07", x"FC43", x"FD03", x"FF61", x"0238", x"03E2", x"04A7", x"04BF", x"03AF", x"0351", x"0549", x"0873", x"0B86", x"0EAC", x"10C5", x"10BE", x"0FD1", x"0E85", x"0C34", x"09C7", x"08CA", x"08D6", x"09D1", x"0C16", x"0E4C", x"0F25", x"0F41", x"0EAE", x"0D46", x"0C7A", x"0CF0", x"0D8B", x"0E46", x"0F63", x"0FA7", x"0F31", x"0F43", x"0F80", x"0F4A", x"0FD7", x"1142", x"126C", x"13ED", x"15B0", x"1628", x"1594", x"1546", x"1525", x"1577", x"177C", x"19CD", x"1AAD", x"1A85", x"1948", x"1689", x"1475", x"145D", x"14CD", x"1585", x"16DE", x"1723", x"15D0", x"1488", x"1300", x"1093", x"0F25", x"0F66", x"100D", x"1174", x"136E", x"13AE", x"11F3", x"0FCA", x"0D24", x"0A6E", x"0988", x"09C4", x"0972", x"092F", x"08BC", x"071D", x"058A", x"050B", x"0484", x"041D", x"04DF", x"05AF", x"0690", x"0891", x"0ABA", x"0C11", x"0DA9", x"0F34", x"0FFC", x"119D", x"1467", x"1609", x"1686", x"1630", x"1379", x"0F6F", x"0D36", x"0C62", x"0B92", x"0C02", x"0CB7", x"0BB4", x"0AC2", x"0B5A", x"0B8C", x"0B73", x"0C99", x"0D8E", x"0DC0", x"0EDB", x"0FC7", x"0E5D", x"0B88", x"07CC", x"027C", x"FD91", x"FAC9", x"F90E", x"F800", x"F82F", x"F83E", x"F785", x"F76F", x"F7AC", x"F77E", x"F803", x"F936", x"FA10", x"FB67", x"FD7E", x"FEF1", x"FFFF", x"018E", x"0284", x"0355", x"059A", x"0860", x"0A1C", x"0B64", x"0BA2", x"09C3", x"0822", x"08D0", x"0AAE", x"0D54", x"1101", x"13AA", x"1430", x"142D", x"13D0", x"1222", x"1057", x"0F3A", x"0E23", x"0D75", x"0DE4", x"0E0E", x"0D20", x"0B90", x"095A", x"06B8", x"0551", x"058E", x"06CF", x"08DC", x"0AF3", x"0BAD", x"0B13", x"09B6", x"078A", x"0559", x"0424", x"0399", x"0356", x"03C2", x"0432", x"03F7", x"042B", x"0502", x"0617", x"086D", x"0C89", x"10F6", x"1495", x"1788", x"186B", x"1720", x"163C", x"1700", x"1897", x"1B07", x"1DF1", x"1F00", x"1DC3", x"1BA6", x"187D", x"1414", x"1038", x"0DB0", x"0BD0", x"0B40", x"0C27", x"0CCA", x"0CA6", x"0C83", x"0BF9", x"0B17", x"0B42", x"0C4A", x"0CEE", x"0D8E", x"0DF2", x"0D07", x"0B79", x"0A2D", x"0861", x"063C", x"04D9", x"03F0", x"034B", x"0409", x"0595", x"06E3", x"08B0", x"0B1C", x"0D66", x"10A2", x"1553", x"197C", x"1C4A", x"1DE5", x"1CEC", x"19B2", x"174A", x"164C", x"1575", x"1583", x"15F5", x"1473", x"11A4", x"0F3F", x"0BF1", x"07C0", x"04DF", x"0344", x"0240", x"0350", x"05EB", x"077B", x"0839", x"08C7", x"0818", x"0736", x"07F3", x"0934", x"09F4", x"0AED", x"0B0F", x"0962", x"0795", x"0632", x"042A", x"02A8", x"0255", x"0257", x"030E", x"0532", x"071D", x"0846", x"09B7", x"0AA0", x"0B05", x"0CA2", x"0EC6", x"0FD4", x"1076", x"1036", x"0D89", x"0A95", x"09E6", x"0A23", x"0B25", x"0D6D", x"0E72", x"0CC3", x"0B14", x"09F9", x"0815", x"06D8", x"06C7", x"05EB", x"04F3", x"05AE", x"065A", x"05DF", x"0539", x"033B", x"FF37", x"FB8C", x"F94F", x"F78B", x"F736", x"F869", x"F907", x"F938", x"FA14", x"FA66", x"FA1F", x"FA9F", x"FB24", x"FB25", x"FBFA", x"FCEB", x"FC6E", x"FB8F", x"FA87", x"F847", x"F696", x"F70E", x"F829", x"F99A", x"FBF6", x"FCD7", x"FB1F", x"F9EF", x"FA74", x"FBCD", x"FF42", x"044F", x"0735", x"07A7", x"07A4", x"0670", x"038E", x"0134", x"FF48", x"FCA2", x"FAE8", x"FABF", x"FA1F", x"F87C", x"F6B5", x"F410", x"F12C", x"EFBC", x"F005", x"F125", x"F36B", x"F612", x"F7DD", x"F8D2", x"F8F8", x"F7F4", x"F6B3", x"F5DE", x"F4FB", x"F460", x"F43B", x"F394", x"F285", x"F209", x"F190", x"F0D1", x"F15B", x"F30A", x"F4BF", x"F6B8", x"F88C", x"F7F7", x"F59E", x"F417", x"F3DF", x"F4FD", x"F856", x"FC1E", x"FD7D", x"FCF3", x"FB9B", x"F8DE", x"F582", x"F377", x"F244", x"F19B", x"F299", x"F482", x"F551", x"F517", x"F432", x"F245", x"F074", x"F018", x"F0BE", x"F22C", x"F4B5", x"F755", x"F920", x"FA9B", x"FB5B", x"FB2C", x"FB64", x"FC36", x"FCB7", x"FD90", x"FEF3", x"FF8C", x"FF87", x"0030", x"005C", x"0029", x"01A7", x"0470", x"0662", x"07C1", x"07DF", x"04BF", x"0008", x"FD23", x"FB85", x"FAC7", x"FBB6", x"FC71", x"FAD0", x"F8B3", x"F712", x"F4A9", x"F25B", x"F190", x"F0D1", x"F044", x"F183", x"F35A", x"F43F", x"F50F", x"F57A", x"F451", x"F346", x"F34F", x"F357", x"F3A0", x"F4D2", x"F552", x"F4C5", x"F450", x"F357", x"F1AC", x"F0C3", x"F087", x"F048", x"F134", x"F327", x"F4B8", x"F683", x"F8BF", x"F9FE", x"FB1D", x"FDB5", x"005F", x"0210", x"0355", x"0245", x"FDC6", x"F8F8", x"F5AB", x"F372", x"F363", x"F58A", x"F6B5", x"F65B", x"F667", x"F5F1", x"F4DA", x"F508", x"F5A3", x"F50D", x"F4D4", x"F576", x"F4F4", x"F3EE", x"F2F8", x"EFF3", x"EB33", x"E74D", x"E3F1", x"E0AA", x"DF2F", x"DEA4", x"DD47", x"DC21", x"DBE6", x"DAF9", x"DA20", x"DA4F", x"DA61", x"DAC5", x"DCE3", x"DFA7", x"E266", x"E624", x"E971", x"EAF6", x"EC7C", x"EE7D", x"EFC5", x"F194", x"F42E", x"F484", x"F2CA", x"F1CB", x"F19A", x"F23B", x"F592", x"F9F8", x"FC09", x"FC91", x"FCA8", x"FB24", x"F91F", x"F866", x"F7AC", x"F643", x"F5E2", x"F5D2", x"F4BA", x"F392", x"F268", x"F019", x"EDE9", x"ED2B", x"ED16", x"ED93", x"EF08", x"EFFD", x"EF97", x"EEA1", x"ED04", x"EAD6", x"E991", x"E972", x"EA1F", x"EBFB", x"EE77", x"F03B", x"F1FA", x"F414", x"F564", x"F675", x"F8B7", x"FB0F", x"FD37", x"005E", x"02E7", x"0259", x"005D", x"FED8", x"FD78", x"FD93", x"0051", x"02C1", x"02CD", x"01D1", x"FFEA", x"FC52", x"F8B5", x"F60C", x"F31C", x"F085", x"EFA9", x"EF85", x"EF58", x"EFEF", x"F043", x"EF71", x"EE76", x"ED96", x"EC3F", x"EB76", x"EBCC", x"EC08", x"EC0D", x"EC57", x"EBDB", x"EA95", x"E9D0", x"E941", x"E8AE", x"E92D", x"EA81", x"EB9E", x"ED53", x"EFAF", x"F17D", x"F381", x"F6E7", x"FA75", x"FDC1", x"015F", x"037A", x"0289", x"00DA", x"FFDB", x"FF0F", x"FFA6", x"01AF", x"0223", x"0003", x"FD0C", x"F952", x"F4DA", x"F1D8", x"F091", x"EFBC", x"F018", x"F1FA", x"F3A9", x"F502", x"F690", x"F747", x"F70B", x"F735", x"F754", x"F6E1", x"F6FB", x"F735", x"F66E", x"F595", x"F50D", x"F3FE", x"F303", x"F2F6", x"F2A3", x"F23A", x"F30E", x"F466", x"F5D2", x"F84A", x"FAC9", x"FBF3", x"FD5E", x"FF8E", x"016D", x"03DA", x"06EE", x"07B4", x"05CB", x"0354", x"0068", x"FD9F", x"FD77", x"FF31", x"FFD3", x"0004", x"0062", x"FF64", x"FDF2", x"FDC6", x"FD1C", x"FB51", x"FA86", x"FA5C", x"F9A7", x"F9AF", x"FA05", x"F873", x"F5CD", x"F392", x"F0DA", x"EE4E", x"ED8F", x"ED9C", x"ED9C", x"EEB4", x"F02A", x"F0B5", x"F101", x"F126", x"F029", x"EF31", x"EF27", x"EF42", x"EFFC", x"F1F9", x"F386", x"F475", x"F615", x"F7F4", x"F9B5", x"FCDF", x"004C", x"0189", x"016B", x"0123", x"0026", x"001C", x"02A8", x"056B", x"0693", x"0705", x"0633", x"03A2", x"01A0", x"00BE", x"FF55", x"FDCF", x"FD2C", x"FC0E", x"FABC", x"FA5F", x"F9D2", x"F80D", x"F697", x"F57D", x"F45B", x"F469", x"F5E8", x"F75B", x"F8A6", x"F9CD", x"F981", x"F7F6", x"F657", x"F455", x"F25C", x"F19A", x"F135", x"F098", x"F102", x"F1F9", x"F221", x"F27B", x"F3CF", x"F4A8", x"F5E8", x"F8AE", x"FA7C", x"F990", x"F7C5", x"F592", x"F314", x"F2E6", x"F5C2", x"F8B4", x"FABC", x"FC88", x"FCC7", x"FB68", x"FA7D", x"F9C8", x"F81D", x"F69F", x"F5D2", x"F49C", x"F3BF", x"F415", x"F442", x"F3F9", x"F452", x"F4D0", x"F4E4", x"F590", x"F6CB", x"F7B2", x"F8DA", x"FA7E", x"FBB4", x"FC5A", x"FCDB", x"FD05", x"FD5B", x"FE94", x"001A", x"01DE", x"0453", x"0694", x"0844", x"0A38", x"0C35", x"0D85", x"0F48", x"1171", x"11AC", x"0F89", x"0C6D", x"085C", x"0481", x"0357", x"0475", x"057A", x"062A", x"0639", x"046B", x"0189", x"FF2E", x"FCDF", x"FAA1", x"F990", x"F915", x"F87D", x"F89E", x"F933", x"F8F8", x"F879", x"F82A", x"F714", x"F5AC", x"F506", x"F426", x"F2C1", x"F1F4", x"F16A", x"F06C", x"EFBB", x"EF3E", x"EE6F", x"EE4D", x"EF84", x"F14C", x"F412", x"F809", x"FB95", x"FE56", x"012E", x"030E", x"03C4", x"0537", x"06B7", x"05FB", x"03B6", x"0155", x"FE42", x"FC42", x"FDC6", x"00B8", x"029D", x"0423", x"0500", x"03EC", x"0288", x"01F3", x"00C3", x"FF15", x"FE62", x"FE06", x"FD63", x"FD76", x"FD78", x"FC3B", x"FA73", x"F887", x"F5C7", x"F342", x"F1CB", x"F0A8", x"EFD7", x"EFF4", x"F001", x"EF78", x"EED9", x"EDEF", x"ECED", x"ECEA", x"EDF6", x"EF93", x"F1F9", x"F489", x"F62C", x"F776", x"F8D9", x"F974", x"FA6C", x"FD12", x"FF96", x"00AC", x"0133", x"00CD", x"FF5C", x"FFB8", x"02D3", x"0648", x"0911", x"0B7D", x"0C20", x"0B01", x"0A1E", x"098A", x"0864", x"07B3", x"079B", x"0725", x"06CB", x"06D6", x"065F", x"058C", x"04F3", x"039C", x"01A2", x"002F", x"FEDD", x"FD46", x"FC71", x"FC11", x"FB11", x"FA60", x"FA77", x"FA2E", x"FA22", x"FB30", x"FC64", x"FDC5", x"0047", x"02F8", x"04D0", x"06D9", x"090B", x"0A86", x"0CCD", x"1052", x"12D0", x"139E", x"13C0", x"12B4", x"1153", x"1242", x"157B", x"1880", x"1AE0", x"1C50", x"1B6E", x"18C3", x"1643", x"13B0", x"110C", x"0F6E", x"0EBF", x"0E19", x"0DBF", x"0DAD", x"0D53", x"0D09", x"0D1C", x"0CCD", x"0C2D", x"0B9A", x"0ACE", x"0A07", x"09F2", x"0A43", x"0A6C", x"0AC1", x"0AE2", x"0A6B", x"0A21", x"0A67", x"0B12", x"0CA3", x"0F29", x"11AD", x"1417", x"16CB", x"191F", x"1B3B", x"1E25", x"2108", x"226B", x"2262", x"2107", x"1DE5", x"1AD9", x"19B7", x"19B6", x"19DD", x"1A55", x"1A1B", x"1869", x"1697", x"157C", x"1470", x"13DE", x"144D", x"14C4", x"14FB", x"1598", x"160F", x"15C9", x"156D", x"14DF", x"1386", x"1204", x"10D8", x"0F86", x"0E76", x"0E5E", x"0EAB", x"0F1C", x"0FE1", x"106A", x"1086", x"110C", x"1229", x"138F", x"15DB", x"18A8", x"1AE7", x"1CDB", x"1EEA", x"2042", x"2178", x"23A6", x"2547", x"24D2", x"22AF", x"1F0E", x"19FB", x"1601", x"1529", x"15F5", x"1776", x"19BD", x"1B7D", x"1BB1", x"1BA0", x"1BB0", x"1B1A", x"1A83", x"1AC0", x"1AFE", x"1B18", x"1B76", x"1BA6", x"1B32", x"1AC1", x"1A32", x"1947", x"184E", x"177A", x"1674", x"15B7", x"1549", x"14B8", x"13E3", x"12A9", x"10A3", x"0E99", x"0D43", x"0C68", x"0C50", x"0D86", x"0EF6", x"0FE0", x"110B", x"11C4", x"116C", x"118E", x"131D", x"1438", x"1428", x"1391", x"11A6", x"0EE3", x"0E27", x"0FFA", x"1286", x"1532", x"17F2", x"1942", x"1923", x"18EE", x"1894", x"17EA", x"17AE", x"17C2", x"1748", x"1645", x"14D2", x"12D4", x"1129", x"1012", x"0F0B", x"0E41", x"0DF2", x"0D4F", x"0C77", x"0BE8", x"0B29", x"09C9", x"08AD", x"0790", x"05E9", x"04BE", x"047B", x"049D", x"059F", x"07C2", x"09C9", x"0B3C", x"0CB4", x"0DAC", x"0DEA", x"0EFC", x"10AA", x"114C", x"108E", x"0EC7", x"0B94", x"0845", x"072D", x"081D", x"09E4", x"0C1C", x"0E19", x"0EA8", x"0DD7", x"0C47", x"0A38", x"083D", x"0712", x"06AA", x"06DD", x"07A7", x"08D0", x"0ACB", x"0DE8", x"1121", x"13BB", x"15D6", x"171B", x"1708", x"167B", x"15F9", x"151F", x"1454", x"144E", x"144A", x"13B8", x"133E", x"1325", x"1369", x"14BA", x"16FF", x"193D", x"1B5A", x"1D51", x"1EBB", x"1FCD", x"2141", x"2239", x"21D4", x"203C", x"1D25", x"18BA", x"14D8", x"1308", x"12AD", x"1326", x"1424", x"1432", x"1292", x"101D", x"0D5F", x"0A4F", x"07E7", x"06B4", x"0641", x"064A", x"0710", x"07D8", x"0882", x"0950", x"09E9", x"09FB", x"0A0C", x"0A2D", x"09C7", x"0943", x"091B", x"08F8", x"08EF", x"0957", x"0990", x"0955", x"095C", x"0A3A", x"0BD3", x"0E21", x"1087", x"126A", x"13AD", x"1482", x"14DC", x"157F", x"169B", x"1768", x"1775", x"169E", x"13E6", x"0FDF", x"0CBA", x"0B95", x"0BBD", x"0D51", x"0F60", x"1022", x"0F4E", x"0E3A", x"0CDA", x"0B19", x"0A0F", x"09EA", x"09DF", x"0A0C", x"0A93", x"0AA1", x"0A21", x"0985", x"0865", x"06A7", x"0482", x"01B9", x"FE4C", x"FAF4", x"F7E4", x"F534", x"F361", x"F246", x"F13E", x"F0AC", x"F088", x"F04C", x"F025", x"F087", x"F09B", x"F0A3", x"F156", x"F224", x"F2D2", x"F4B4", x"F7A3", x"FA20", x"FC21", x"FD4B", x"FC6B", x"FA9E", x"FAA7", x"FC6E", x"FEFF", x"024E", x"0555", x"0639", x"059F", x"04CC", x"0341", x"013A", x"FFE4", x"FF1F", x"FE21", x"FCF3", x"FB7D", x"F985", x"F7B6", x"F6BC", x"F6A2", x"F73A", x"F803", x"F89E", x"F946", x"FA36", x"FB0E", x"FBFE", x"FD13", x"FD74", x"FD23", x"FCCA", x"FC2A", x"FB44", x"FB18", x"FBB2", x"FC69", x"FD78", x"FEC3", x"FF48", x"FF4A", x"FFED", x"00BE", x"0138", x"0194", x"0130", x"FF88", x"FDED", x"FDB6", x"FE85", x"0012", x"0234", x"03A9", x"03AA", x"027F", x"0062", x"FD7C", x"FA73", x"F7DE", x"F583", x"F35C", x"F12B", x"EEE3", x"ED2C", x"EC5C", x"EC0F", x"EC3A", x"ECC1", x"ECEC", x"EC85", x"EC4D", x"EC2B", x"EBF8", x"EC68", x"EDDE", x"EF5C", x"F0B3", x"F204", x"F31D", x"F400", x"F5B8", x"F82E", x"FAC9", x"FD6A", x"FFD9", x"01A4", x"0310", x"0489", x"0568", x"053B", x"03EA", x"011A", x"FD11", x"F97D", x"F752", x"F6A9", x"F77C", x"F97B", x"FB27", x"FC04", x"FC49", x"FBE9", x"FAD6", x"F9E9", x"F955", x"F8C4", x"F85A", x"F826", x"F7A8", x"F6E8", x"F650", x"F574", x"F465", x"F383", x"F2A5", x"F15C", x"F03B", x"EFA4", x"EF69", x"EFD0", x"F0E5", x"F1E8", x"F26B", x"F2EA", x"F3D8", x"F55B", x"F797", x"FA43", x"FD2B", x"FFDB", x"01EE", x"0339", x"0413", x"042B", x"0370", x"0259", x"0089", x"FCEE", x"F897", x"F565", x"F3C6", x"F3FF", x"F6B7", x"FA1C", x"FC21", x"FCE7", x"FD2F", x"FC40", x"FAA7", x"F9A9", x"F8BB", x"F775", x"F6BA", x"F661", x"F57A", x"F471", x"F3C3", x"F2EC", x"F1ED", x"F10D", x"EF74", x"ECD8", x"E9EA", x"E74A", x"E546", x"E48B", x"E4E5", x"E5CD", x"E72B", x"E8C1", x"EA87", x"ECB6", x"EF23", x"F168", x"F3FC", x"F680", x"F7CA", x"F838", x"F8AB", x"F8AD", x"F875", x"F8EB", x"F8B5", x"F675", x"F3C2", x"F254", x"F1C3", x"F2A7", x"F56F", x"F846", x"F999", x"FA7A", x"FAF8", x"FA2B", x"F8C4", x"F7C9", x"F6F0", x"F5F0", x"F52E", x"F441", x"F2CD", x"F17E", x"F0F1", x"F136", x"F1C8", x"F1D3", x"F0F5", x"EF5C", x"ED12", x"EABF", x"E917", x"E7FA", x"E6EA", x"E686", x"E6AD", x"E696", x"E6CF", x"E7D8", x"E927", x"EAD4", x"EDB1", x"F078", x"F1F4", x"F2EC", x"F3C3", x"F3F8", x"F44D", x"F529", x"F4E2", x"F2E1", x"F0C2", x"EF3F", x"EDF8", x"EDCE", x"EE9D", x"EF07", x"EE91", x"EDF3", x"ECD9", x"EB01", x"E927", x"E81F", x"E7D2", x"E85E", x"E9A6", x"EB7A", x"ED99", x"F016", x"F2D9", x"F58A", x"F78E", x"F84C", x"F7F4", x"F6D3", x"F528", x"F3A0", x"F2F0", x"F313", x"F3A7", x"F4AA", x"F5A8", x"F69C", x"F7F0", x"FA26", x"FCF9", x"002B", x"035C", x"05A5", x"06C0", x"073E", x"0763", x"0740", x"0739", x"06F1", x"055E", x"0299", x"FFB6", x"FD2B", x"FB58", x"FAEE", x"FB61", x"FB8B", x"FB25", x"FA6D", x"F8FD", x"F708", x"F58A", x"F4A2", x"F415", x"F402", x"F425", x"F3E6", x"F37D", x"F32A", x"F2B3", x"F22A", x"F193", x"F08F", x"EED9", x"ECF0", x"EB03", x"E965", x"E8C4", x"E8FC", x"E963", x"E985", x"E964", x"E920", x"E96F", x"EABE", x"ECEE", x"EFEC", x"F356", x"F632", x"F889", x"FAE1", x"FD01", x"FF21", x"01EC", x"041D", x"03DB", x"01EC", x"FF90", x"FD06", x"FBBC", x"FCDD", x"FE93", x"FEFF", x"FED6", x"FDE5", x"FB46", x"F828", x"F5C8", x"F384", x"F197", x"F12D", x"F169", x"F13A", x"F125", x"F14E", x"F136", x"F14C", x"F1B1", x"F16D", x"F023", x"EE42", x"EC27", x"EA70", x"E997", x"E960", x"E954", x"E8F0", x"E7D9", x"E652", x"E4F8", x"E37B", x"E264", x"E273", x"E30A", x"E355", x"E41B", x"E55A", x"E67F", x"E8CD", x"ECCB", x"F038", x"F1F0", x"F323", x"F3EB", x"F47A", x"F6BD", x"FAC3", x"FE2A", x"006D", x"022C", x"028C", x"0145", x"FF8C", x"FD96", x"FAE7", x"F852", x"F627", x"F3DD", x"F190", x"EFF4", x"EF66", x"F03A", x"F223", x"F44F", x"F61A", x"F71D", x"F6F9", x"F64D", x"F5B0", x"F4C9", x"F3BE", x"F33E", x"F2D7", x"F217", x"F1F7", x"F26D", x"F2CE", x"F3ED", x"F61E", x"F7DF", x"F8AE", x"F960", x"F9CF", x"F9F2", x"FB45", x"FD71", x"FE52", x"FDC3", x"FCF8", x"FC03", x"FBC2", x"FD82", x"009E", x"0330", x"0520", x"068C", x"06A6", x"0570", x"03D3", x"0207", x"FFDA", x"FDFA", x"FC9F", x"FB69", x"FA4A", x"FA28", x"FB3E", x"FD2F", x"FF81", x"018F", x"0285", x"022E", x"0146", x"00B5", x"009F", x"0112", x"0206", x"02E8", x"0340", x"036C", x"03EA", x"04BC", x"05E6", x"07C5", x"098D", x"0A34", x"09AF", x"087D", x"06DA", x"05AA", x"05F7", x"06E0", x"06FC", x"065C", x"0580", x"04B0", x"04F5", x"0775", x"0AF0", x"0E05", x"1085", x"11F0", x"1177", x"0FD8", x"0E19", x"0BE8", x"0954", x"073A", x"0520", x"025D", x"FFB2", x"FD5A", x"FB16", x"F95B", x"F885", x"F7C9", x"F6BF", x"F5B2", x"F4A7", x"F425", x"F4D9", x"F6C2", x"F928", x"FBD4", x"FE11", x"FFE6", x"01F3", x"0447", x"06B1", x"0974", x"0BE4", x"0C72", x"0B5A", x"0964", x"068E", x"03F5", x"02FD", x"0237", x"000C", x"FD99", x"FB68", x"F99A", x"F9F5", x"FD53", x"014E", x"04A5", x"07C4", x"0961", x"08E2", x"07EB", x"0709", x"058B", x"048E", x"04DB", x"051E", x"0518", x"0548", x"04E7", x"03C2", x"02C3", x"01D3", x"0025", x"FDF5", x"FB56", x"F85D", x"F5FA", x"F4B3", x"F443", x"F4B4", x"F5A1", x"F68C", x"F7CB", x"F978", x"FA8A", x"FB7B", x"FCCC", x"FD5D", x"FCCF", x"FC45", x"FB5D", x"FA19", x"FA8F", x"FC9C", x"FDBA", x"FD44", x"FC17", x"F98B", x"F720", x"F77D", x"F9D8", x"FC37", x"FEBD", x"0102", x"0199", x"0193", x"01F6", x"01DA", x"0115", x"00A4", x"FFE4", x"FE69", x"FD4F", x"FCB9", x"FC33", x"FC48", x"FCF9", x"FD2F", x"FCB2", x"FB9A", x"F98D", x"F745", x"F5AE", x"F4C7", x"F49C", x"F551", x"F61A", x"F6EA", x"F858", x"F9D6", x"FAEF", x"FC81", x"FE0F", x"FE83", x"FE4C", x"FDFA", x"FCE0", x"FC02", x"FD11", x"FE9A", x"FEAE", x"FD6C", x"FAD4", x"F6CF", x"F3C7", x"F388", x"F4D2", x"F685", x"F8A4", x"FA52", x"FAA1", x"FAC6", x"FB4A", x"FBCD", x"FC9A", x"FE4F", x"0028", x"019C", x"0313", x"04B2", x"0670", x"0889", x"0AD5", x"0C8F", x"0CFD", x"0C2F", x"0A7C", x"0892", x"06F7", x"061A", x"0628", x"06B7", x"077D", x"0910", x"0B5C", x"0DF0", x"10EB", x"1490", x"17C1", x"19B3", x"1AE1", x"1B17", x"1A05", x"1955", x"1A12", x"1AAA", x"19E3", x"17E9", x"1444", x"0F19", x"0B0C", x"0970", x"08C0", x"0877", x"08DB", x"08A4", x"0736", x"0610", x"053B", x"03E8", x"02E3", x"0302", x"031C", x"02EA", x"0321", x"031F", x"02B2", x"02C8", x"036E", x"03CE", x"03F8", x"03F7", x"0354", x"0276", x"01E8", x"0166", x"012C", x"0154", x"0183", x"0223", x"03AD", x"05B8", x"0847", x"0BB4", x"0EE8", x"10E7", x"12AC", x"142B", x"1509", x"16C5", x"19AB", x"1B5F", x"1B20", x"199F", x"1681", x"12A5", x"1121", x"11FF", x"1339", x"14A7", x"15DC", x"14F1", x"12A4", x"10A7", x"0E44", x"0B52", x"097B", x"086E", x"0758", x"0722", x"07B2", x"07C1", x"07BB", x"083E", x"0831", x"07A3", x"070B", x"05B7", x"03B5", x"01F7", x"0030", x"FE3E", x"FD13", x"FC51", x"FB87", x"FBAC", x"FC78", x"FCC2", x"FD5D", x"FE78", x"FE7B", x"FDED", x"FE26", x"FE83", x"FF7F", x"032E", x"082C", x"0BD3", x"0E37", x"0EDF", x"0CEE", x"0B14", x"0C04", x"0E84", x"1179", x"14FD", x"16C8", x"15A6", x"13B5", x"11A8", x"0E85", x"0B7C", x"0977", x"072A", x"050A", x"047C", x"04AC", x"052B", x"0710", x"0A12", x"0D06", x"0FE3", x"1212", x"1284", x"11A0", x"101F", x"0E03", x"0C3C", x"0B35", x"0A99", x"0ACC", x"0C0F", x"0D00", x"0D64", x"0E0E", x"0E27", x"0D4F", x"0CD2", x"0CAD", x"0BE0", x"0C53", x"0EF6", x"11F3", x"143F", x"1611", x"15C3", x"1384", x"1265", x"1363", x"153F", x"17DA", x"1A8C", x"1AD0", x"18CC", x"1636", x"12D8", x"0E9F", x"0B10", x"081E", x"0500", x"0277", x"0134", x"0048", x"0009", x"012F", x"0350", x"05B6", x"0854", x"0A50", x"0B2C", x"0B52", x"0AFE", x"0AA0", x"0AE4", x"0BD9", x"0D75", x"1052", x"13DC", x"1685", x"1863", x"19A8", x"196B", x"1811", x"1709", x"15D1", x"140E", x"13C7", x"1561", x"16C9", x"1785", x"17B6", x"162B", x"1384", x"12C3", x"13ED", x"157E", x"1781", x"1988", x"19E9", x"1931", x"18E8", x"1867", x"175B", x"16DD", x"165E", x"14E3", x"130C", x"113C", x"0EB2", x"0C0B", x"0A3E", x"08B0", x"0760", x"0699", x"05DE", x"04D6", x"0410", x"039A", x"0372", x"041A", x"056F", x"0742", x"0A33", x"0DC0", x"10D8", x"13AD", x"1628", x"16F3", x"16A7", x"1630", x"14CE", x"12C8", x"1284", x"1374", x"13D7", x"13EA", x"1376", x"1131", x"0F29", x"1006", x"129F", x"15C5", x"1975", x"1BE0", x"1B6F", x"19EA", x"1829", x"155E", x"12CC", x"1148", x"0F63", x"0D39", x"0BE7", x"0A63", x"0836", x"06BB", x"05A6", x"0417", x"0369", x"0392", x"02FB", x"020E", x"0170", x"0070", x"FFC9", x"00D4", x"0299", x"049A", x"076C", x"09F9", x"0B24", x"0C04", x"0C33", x"0ACE", x"094B", x"0845", x"06A6", x"05C0", x"074B", x"098F", x"0B48", x"0CE4", x"0C97", x"099C", x"075D", x"07A4", x"095E", x"0CDE", x"11DE", x"158D", x"1766", x"1923", x"1A06", x"1978", x"18F0", x"1827", x"15E0", x"135D", x"111C", x"0E23", x"0B09", x"08FC", x"0704", x"0535", x"0476", x"03B0", x"021F", x"0042", x"FE1B", x"FB6C", x"F9CF", x"F9B4", x"FAC5", x"FD69", x"011E", x"03D7", x"058D", x"0664", x"058C", x"03FD", x"0396", x"034E", x"028C", x"0332", x"04ED", x"05D3", x"065D", x"0633", x"02E9", x"FDB4", x"FA31", x"F87C", x"F808", x"F999", x"FB99", x"FB73", x"FA74", x"F9FF", x"F926", x"F856", x"F8BF", x"F931", x"F91C", x"F9C4", x"FADD", x"FBBB", x"FD59", x"FFED", x"024E", x"04B4", x"0704", x"0801", x"0762", x"05DD", x"031B", x"FFA9", x"FD24", x"FBCD", x"FBE4", x"FE1D", x"01A0", x"04CD", x"07C2", x"0A1F", x"0ACD", x"0AC0", x"0ADB", x"09F5", x"086B", x"081E", x"0892", x"0862", x"0836", x"0747", x"03CC", x"FF8E", x"FD11", x"FBD4", x"FB6E", x"FC95", x"FDC2", x"FD9C", x"FD7B", x"FE1B", x"FE7E", x"FF08", x"0017", x"0029", x"FEEF", x"FD0B", x"FA3C", x"F6A6", x"F3DB", x"F1EE", x"F068", x"EFC5", x"EF7D", x"EE43", x"EC60", x"EA1C", x"E719", x"E44D", x"E320", x"E32B", x"E49B", x"E7E1", x"EB8B", x"EE82", x"F1A0", x"F46C", x"F629", x"F80C", x"FA4D", x"FB36", x"FBEF", x"FE08", x"0053", x"01EF", x"03CD", x"041E", x"01BA", x"FF54", x"FEA4", x"FE87", x"FF74", x"01A8", x"024F", x"00FC", x"FF90", x"FDB0", x"FB0B", x"F965", x"F896", x"F724", x"F658", x"F6B8", x"F69A", x"F644", x"F681", x"F5D3", x"F430", x"F354", x"F299", x"F0B8", x"EEB6", x"EC57", x"E8A4", x"E549", x"E345", x"E1C1", x"E12A", x"E1E8", x"E25B", x"E22C", x"E276", x"E22E", x"E141", x"E155", x"E1BE", x"E150", x"E22E", x"E50B", x"E823", x"EBC3", x"EFEC", x"F1BD", x"F13F", x"F1A1", x"F31E", x"F523", x"F8FA", x"FD46", x"FF46", x"FFD3", x"0041", x"FF51", x"FDE3", x"FD4A", x"FBF5", x"F974", x"F7AB", x"F65F", x"F4C5", x"F489", x"F56F", x"F5E8", x"F6B5", x"F86F", x"F95C", x"F92D", x"F88E", x"F66F", x"F312", x"F092", x"EF0E", x"EEA5", x"F086", x"F38D", x"F598", x"F703", x"F77C", x"F5BF", x"F3BE", x"F330", x"F259", x"F1A3", x"F35A", x"F673", x"F96E", x"FD38", x"002D", x"FF38", x"FC53", x"FA8B", x"F98B", x"F9FB", x"FCEB", x"FFA9", x"001C", x"FFB2", x"FEA3", x"FC32", x"FA04", x"F8DD", x"F72C", x"F586", x"F502", x"F495", x"F45A", x"F5AD", x"F790", x"F910", x"FB16", x"FD20", x"FDAC", x"FD53", x"FC29", x"F95D", x"F612", x"F3EB", x"F28A", x"F28D", x"F497", x"F6BC", x"F7DA", x"F888", x"F817", x"F60A", x"F49C", x"F419", x"F2DA", x"F209", x"F357", x"F54D", x"F7AB", x"FB63", x"FE2B", x"FE25", x"FD9D", x"FE06", x"FE71", x"FFCC", x"0269", x"03EA", x"03FB", x"045D", x"04B9", x"04E1", x"0604", x"0750", x"06F4", x"059A", x"0357", x"FF55", x"FB1E", x"F830", x"F590", x"F392", x"F36E", x"F3E5", x"F3BE", x"F3CA", x"F32B", x"F0DB", x"EE9E", x"EDD7", x"EDCC", x"EF56", x"F2A9", x"F598", x"F775", x"F918", x"F964", x"F812", x"F70D", x"F5D6", x"F333", x"F160", x"F14E", x"F193", x"F2C8", x"F567", x"F680", x"F582", x"F542", x"F607", x"F732", x"FA4A", x"FE60", x"006E", x"0115", x"0192", x"00D1", x"FF82", x"FF2B", x"FE3D", x"FC1C", x"FA86", x"F941", x"F78B", x"F714", x"F7A4", x"F71C", x"F669", x"F67F", x"F5E1", x"F4C8", x"F475", x"F369", x"F12D", x"EFE5", x"EF90", x"EF48", x"F055", x"F229", x"F2BF", x"F2E0", x"F335", x"F258", x"F137", x"F143", x"F092", x"EEDC", x"EE79", x"EEE4", x"EF38", x"F142", x"F3E9", x"F3A7", x"F1B5", x"F08A", x"EF6C", x"EF7E", x"F2A9", x"F63C", x"F7BC", x"F910", x"FA3F", x"FA46", x"FACC", x"FC4E", x"FC4E", x"FB1F", x"FA38", x"F85D", x"F5E6", x"F4A1", x"F38F", x"F1B2", x"F0EE", x"F103", x"F08D", x"F097", x"F122", x"F00C", x"EE2C", x"ED45", x"EC86", x"EC8E", x"EED4", x"F18C", x"F30D", x"F43D", x"F43C", x"F1EB", x"EF94", x"EDD6", x"EB25", x"E8E1", x"E8B9", x"E938", x"EA7D", x"EDC4", x"F01E", x"EF1B", x"ED09", x"EB25", x"E93A", x"E9C7", x"ED69", x"F0B2", x"F2AC", x"F48B", x"F534", x"F494", x"F4A9", x"F4F8", x"F43B", x"F3D9", x"F411", x"F3E8", x"F4C7", x"F775", x"FA27", x"FCE6", x"0037", x"0254", x"02E1", x"038B", x"0350", x"0130", x"FF3A", x"FE1E", x"FD32", x"FE21", x"019F", x"0505", x"07A5", x"0A3E", x"0B2E", x"0A4C", x"09AB", x"08B0", x"0613", x"03C1", x"026A", x"00AE", x"FFDB", x"004D", x"FF15", x"FB84", x"F816", x"F4C8", x"F1F6", x"F1DB", x"F3A2", x"F44F", x"F482", x"F523", x"F523", x"F569", x"F743", x"F8F4", x"F94D", x"F949", x"F815", x"F538", x"F2C1", x"F12E", x"EF69", x"EE8A", x"EEF7", x"EF09", x"EF16", x"F010", x"F045", x"EF35", x"EECD", x"EF0B", x"EF95", x"F1F5", x"F5DD", x"F937", x"FC67", x"FFAB", x"01A5", x"02BA", x"0410", x"046F", x"03D6", x"0437", x"0529", x"0645", x"0920", x"0CA2", x"0DFC", x"0DAB", x"0CDB", x"0AA8", x"08BC", x"091E", x"09CD", x"090F", x"083D", x"06F5", x"046B", x"02C4", x"0280", x"0187", x"004A", x"FFB9", x"FE84", x"FD26", x"FD8C", x"FE3E", x"FDFA", x"FE09", x"FDDE", x"FC3A", x"FACE", x"FA16", x"F80D", x"F55D", x"F397", x"F1CB", x"F055", x"F0DB", x"F210", x"F2B4", x"F3D4", x"F4E3", x"F47A", x"F427", x"F421", x"F2B9", x"F0EF", x"F053", x"EFA9", x"EFA6", x"F220", x"F4A5", x"F4C1", x"F3EE", x"F2C8", x"F0CF", x"F0CA", x"F406", x"F75E", x"F9C8", x"FC4A", x"FDCB", x"FDFF", x"FF04", x"0050", x"005D", x"0022", x"FFF2", x"FED5", x"FDEB", x"FE48", x"FE4F", x"FE09", x"FE55", x"FE13", x"FD11", x"FCD5", x"FCAD", x"FB76", x"FA5F", x"F9A4", x"F880", x"F84E", x"F9C8", x"FB9C", x"FDEB", x"00C1", x"024F", x"0257", x"0276", x"01E1", x"0060", x"FFF1", x"0093", x"00EF", x"030B", x"06DE", x"08F8", x"087F", x"06F8", x"03DA", x"0032", x"FF5B", x"00B7", x"0181", x"01CA", x"0175", x"FF05", x"FBEC", x"F9F8", x"F82D", x"F69E", x"F634", x"F59D", x"F470", x"F49C", x"F5DC", x"F6E1", x"F8C6", x"FB4F", x"FC66", x"FD36", x"FEE7", x"FFB7", x"FF25", x"FF05", x"FEB3", x"FDFC", x"FED6", x"0165", x"03D7", x"06AC", x"099C", x"0ACB", x"0AB3", x"0A82", x"0932", x"0719", x"0630", x"05D3", x"05C0", x"07E7", x"0B53", x"0CFB", x"0D04", x"0C47", x"0A08", x"07CA", x"07E4", x"08F3", x"093E", x"0993", x"09A2", x"08C4", x"0846", x"08D7", x"0943", x"09B8", x"09F3", x"08AB", x"063D", x"0413", x"01C2", x"FF7B", x"FE5B", x"FD6D", x"FBCE", x"FAC2", x"FA49", x"F8E7", x"F74D", x"F65E", x"F571", x"F517", x"F650", x"F84C", x"FA7C", x"FD55", x"FFC2", x"00E7", x"01D1", x"0239", x"01D1", x"0239", x"03C1", x"04DD", x"06B3", x"0A57", x"0D84", x"0EF6", x"0FF5", x"0FAB", x"0DC7", x"0D72", x"0F7C", x"1157", x"127B", x"134D", x"1208", x"0F39", x"0D44", x"0BE6", x"0A38", x"0966", x"08E5", x"076B", x"068B", x"071E", x"07AD", x"0872", x"0A0F", x"0AE3", x"0AA3", x"0B39", x"0BED", x"0B77", x"0B14", x"0AEE", x"0A17", x"0964", x"09C6", x"0A13", x"0A62", x"0B82", x"0C46", x"0C45", x"0C43", x"0B94", x"09D0", x"089B", x"07FF", x"0751", x"0841", x"0B48", x"0DDF", x"0F26", x"0FCC", x"0ED5", x"0CCA", x"0CD3", x"0EEF", x"10F9", x"12CD", x"147B", x"14B2", x"141D", x"1444", x"1453", x"1397", x"1292", x"10C1", x"0DA6", x"0A6D", x"0764", x"0483", x"0279", x"0147", x"FFD6", x"FE83", x"FD9B", x"FC6A", x"FB52", x"FB35", x"FB51", x"FBB2", x"FD53", x"FFA0", x"01F1", x"04EF", x"07AE", x"087D", x"083C", x"079E", x"059C", x"039C", x"032A", x"0314", x"0346", x"05E7", x"09B9", x"0C1E", x"0D8E", x"0DEE", x"0BDD", x"09B9", x"0A8F", x"0CD8", x"0F1C", x"11BC", x"12F3", x"1171", x"0F5E", x"0DBF", x"0B90", x"099C", x"08CC", x"0785", x"062F", x"064C", x"0701", x"07CA", x"09E7", x"0C49", x"0DAA", x"0F1B", x"10C0", x"110B", x"10BB", x"10A5", x"0F93", x"0E25", x"0E08", x"0E84", x"0EFB", x"108C", x"123B", x"129A", x"12D6", x"131B", x"11EC", x"1034", x"0F17", x"0D75", x"0C16", x"0CDF", x"0E58", x"0EE2", x"0F41", x"0F14", x"0DA5", x"0D1B", x"0EB1", x"1084", x"120F", x"1393", x"13AC", x"129C", x"122B", x"1250", x"1230", x"126E", x"1216", x"0FDB", x"0CBC", x"0970", x"05AB", x"0265", x"008E", x"FEB0", x"FCDD", x"FBE1", x"FAED", x"F9BB", x"F993", x"FA10", x"FA72", x"FBE7", x"FE7A", x"00E2", x"03DF", x"0783", x"09D8", x"0B0A", x"0C47", x"0C77", x"0B91", x"0BBC", x"0C32", x"0C18", x"0D8A", x"10F8", x"13D2", x"1609", x"1803", x"17B5", x"15D5", x"15CF", x"175B", x"18E6", x"1B16", x"1CC8", x"1BE1", x"19CF", x"1892", x"1709", x"1571", x"14D4", x"139B", x"111A", x"0F49", x"0E26", x"0CBC", x"0BF2", x"0BA8", x"0A0C", x"079D", x"0596", x"02EE", x"FFF0", x"FE08", x"FCB3", x"FB8B", x"FB73", x"FBF7", x"FBDF", x"FC05", x"FC8E", x"FC7A", x"FCAE", x"FD8B", x"FDD2", x"FDA1", x"FDDF", x"FD60", x"FC24", x"FC69", x"FE03", x"FF65", x"0119", x"02B5", x"0298", x"0241", x"043B", x"07B1", x"0B95", x"1037", x"1434", x"1609", x"1740", x"1886", x"1914", x"1942", x"1977", x"18A2", x"16B7", x"14D0", x"1294", x"102C", x"0E81", x"0CE9", x"0AA8", x"0892", x"06B8", x"0459", x"029E", x"01DE", x"013B", x"010E", x"0234", x"0370", x"049F", x"06A0", x"0853", x"08C7", x"0924", x"090D", x"077D", x"05FC", x"0531", x"038D", x"025D", x"03BC", x"0622", x"082F", x"0AB3", x"0BBE", x"09BF", x"07E3", x"086F", x"09A1", x"0B71", x"0E51", x"0FAC", x"0EDA", x"0E4C", x"0E00", x"0CC0", x"0BE7", x"0BA3", x"0A87", x"0997", x"09D9", x"0A33", x"0AD4", x"0C90", x"0DB2", x"0DBF", x"0E09", x"0E0F", x"0D07", x"0C96", x"0CA2", x"0BFE", x"0BC5", x"0CE2", x"0D92", x"0E08", x"0F40", x"0FEA", x"0FD0", x"1067", x"10E8", x"1056", x"102B", x"100F", x"0EC6", x"0E51", x"0FD0", x"115A", x"12DA", x"14C7", x"14B2", x"128D", x"11EB", x"1304", x"144A", x"1684", x"18D3", x"18B5", x"1759", x"1707", x"16DA", x"16D8", x"180A", x"18CD", x"17C7", x"164D", x"1419", x"10CB", x"0E0B", x"0C11", x"0935", x"0678", x"049B", x"0239", x"FFD2", x"FEAB", x"FD42", x"FB1F", x"FA3B", x"FA0B", x"F962", x"F987", x"FA49", x"F9F9", x"F9B8", x"FA76", x"FA85", x"FA5C", x"FB0C", x"FAD7", x"F9A5", x"FA19", x"FBE8", x"FDBA", x"00AE", x"03AE", x"03C2", x"0282", x"02D6", x"03B0", x"04F6", x"07C7", x"09C1", x"0906", x"07DB", x"073E", x"061F", x"0595", x"0616", x"05A8", x"0479", x"0403", x"03D7", x"03F1", x"05A1", x"079F", x"0892", x"0932", x"094C", x"07EF", x"0651", x"052C", x"037D", x"01ED", x"0149", x"005E", x"FEE2", x"FDC5", x"FC45", x"FA21", x"F8D4", x"F816", x"F6FF", x"F6B8", x"F6F4", x"F5BF", x"F427", x"F3A3", x"F32C", x"F2F8", x"F43D", x"F4E6", x"F33C", x"F1C9", x"F1E7", x"F2AF", x"F50C", x"F925", x"FBF2", x"FC9C", x"FD39", x"FD8E", x"FD58", x"FDFF", x"FF30", x"FF11", x"FE67", x"FDEC", x"FCC1", x"FB67", x"FAD5", x"F9D3", x"F80D", x"F6B0", x"F563", x"F3BA", x"F2CB", x"F2B7", x"F26F", x"F299", x"F34E", x"F356", x"F2F4", x"F2CE", x"F209", x"F0B6", x"EFCF", x"EE6E", x"EC34", x"EA8C", x"E8E2", x"E629", x"E44F", x"E48B", x"E589", x"E7AA", x"EB25", x"ED13", x"EC89", x"EC50", x"ED38", x"EE57", x"F0E2", x"F44F", x"F5C6", x"F560", x"F4FE", x"F3ED", x"F20B", x"F0F7", x"EFFF", x"EE31", x"ED03", x"ECE8", x"ED2C", x"EE92", x"F199", x"F4B3", x"F7A6", x"FAE1", x"FD1E", x"FE0E", x"FEDD", x"FF5F", x"FF83", x"005C", x"018C", x"021C", x"02D5", x"0381", x"032B", x"028C", x"0208", x"0054", x"FE4A", x"FD39", x"FB56", x"F855", x"F685", x"F586", x"F44C", x"F470", x"F551", x"F3BD", x"F106", x"F021", x"F054", x"F185", x"F515", x"F861", x"F8BE", x"F810", x"F787", x"F61A", x"F55B", x"F631", x"F656", x"F550", x"F4AE", x"F383", x"F192", x"F0B2", x"F08E", x"EFD4", x"EFAF", x"F057", x"F052", x"F047", x"F114", x"F1CE", x"F2D7", x"F53C", x"F7CC", x"F9B7", x"FBA9", x"FCB0", x"FC59", x"FC1B", x"FBF4", x"FB1B", x"FAEC", x"FB71", x"FAA8", x"F961", x"F95C", x"F9C5", x"FAD5", x"FE04", x"0122", x"01CB", x"01C6", x"0224", x"01FC", x"025D", x"03E3", x"0400", x"0208", x"0003", x"FDE5", x"FB76", x"FA06", x"F94A", x"F7A4", x"F587", x"F3A8", x"F19D", x"F02F", x"F04E", x"F134", x"F24F", x"F384", x"F3D5", x"F2FD", x"F1D3", x"F092", x"EF91", x"EFC8", x"F083", x"F0D7", x"F132", x"F14C", x"F03F", x"EF1D", x"EEA8", x"EDB3", x"ECEA", x"EDA3", x"EE39", x"ED55", x"EC5A", x"EB6C", x"E9A4", x"E92F", x"EA9D", x"EB36", x"EA48", x"E9F9", x"EA28", x"EB0D", x"EE93", x"F3EB", x"F7E4", x"FA9C", x"FD09", x"FE38", x"FE5C", x"FF16", x"FF5F", x"FE20", x"FC97", x"FB46", x"F968", x"F789", x"F65F", x"F4E0", x"F2E5", x"F115", x"EF4C", x"ED62", x"EC3F", x"EC4A", x"ED7E", x"EFFB", x"F317", x"F5BB", x"F7C2", x"F905", x"F972", x"F9D5", x"FA89", x"FAD6", x"FAE1", x"FB23", x"FA90", x"F8DB", x"F74A", x"F625", x"F525", x"F55A", x"F677", x"F662", x"F506", x"F404", x"F371", x"F383", x"F553", x"F799", x"F81D", x"F73E", x"F5E7", x"F389", x"F0E2", x"EF55", x"EE38", x"ECD6", x"EC11", x"EBF4", x"EB8B", x"EB83", x"EC80", x"EDFA", x"EFAE", x"F198", x"F31F", x"F3D9", x"F461", x"F552", x"F73C", x"F9E9", x"FC94", x"FEC6", x"0092", x"015B", x"018D", x"022B", x"0294", x"0256", x"02B2", x"0384", x"031E", x"01F4", x"011C", x"FF8F", x"FDFB", x"FE2B", x"FE89", x"FCE6", x"FAEE", x"F9C7", x"F8E8", x"F9FA", x"FDFC", x"019E", x"0331", x"045D", x"04CA", x"03D8", x"039F", x"0454", x"0390", x"01B7", x"0018", x"FDA8", x"FA41", x"F7B5", x"F5AE", x"F355", x"F1B1", x"F0A4", x"EEBE", x"EC48", x"EA0E", x"E83E", x"E7CC", x"E92B", x"EB5A", x"ED83", x"EF51", x"EFE5", x"EFB8", x"EFE2", x"F02A", x"F0C1", x"F2BB", x"F541", x"F6BA", x"F7D9", x"F8F0", x"F932", x"FA01", x"FC72", x"FE86", x"FF16", x"FF9A", x"0010", x"0021", x"0158", x"03A4", x"049E", x"0414", x"034F", x"01E2", x"FFCD", x"FE6F", x"FD9D", x"FC62", x"FB64", x"FB36", x"FB66", x"FBE2", x"FD2A", x"FF05", x"00D3", x"01FC", x"020B", x"00E4", x"FEBE", x"FC75", x"FB7C", x"FBCB", x"FC2C", x"FC34", x"FBF7", x"FA91", x"F880", x"F786", x"F740", x"F6D8", x"F7A1", x"F99F", x"FAA8", x"FA65", x"F9CA", x"F7DB", x"F510", x"F42C", x"F507", x"F528", x"F4CC", x"F4D6", x"F463", x"F46D", x"F6F5", x"FA87", x"FCE9", x"FEB5", x"0065", x"00EF", x"0142", x"0245", x"02CB", x"01FE", x"00ED", x"FF9D", x"FD88", x"FB7F", x"FA12", x"F8B4", x"F770", x"F68C", x"F573", x"F3E3", x"F293", x"F1F9", x"F26F", x"F43B", x"F6BC", x"F8F5", x"FA81", x"FB27", x"FB22", x"FB46", x"FC0D", x"FD04", x"FE3B", x"FF65", x"FF8A", x"FE9C", x"FDD2", x"FD67", x"FD8C", x"FF1A", x"011B", x"019E", x"0099", x"FF5F", x"FDFB", x"FD42", x"FE70", x"0048", x"00C7", x"0042", x"FF12", x"FC85", x"F96C", x"F74B", x"F5B5", x"F476", x"F482", x"F58C", x"F66F", x"F773", x"F906", x"FA90", x"FBFD", x"FD5A", x"FDEB", x"FD38", x"FC08", x"FB38", x"FB62", x"FCAA", x"FE7F", x"0011", x"0092", x"FF9D", x"FDE1", x"FC24", x"FA6A", x"F947", x"F98E", x"FA63", x"FAAC", x"FAD3", x"FAA6", x"F943", x"F837", x"F8E7", x"F97F", x"F931", x"F953", x"F99E", x"F9BA", x"FC12", x"009A", x"041A", x"05F6", x"0745", x"070E", x"05B7", x"05C5", x"0646", x"0524", x"037C", x"01E2", x"FF30", x"FC48", x"FAC7", x"F92F", x"F765", x"F6B1", x"F68C", x"F5B7", x"F51D", x"F4E1", x"F472", x"F4E4", x"F6D1", x"F90E", x"FB0F", x"FC99", x"FCBB", x"FBED", x"FB57", x"FAE5", x"FB18", x"FCE6", x"FF06", x"006A", x"01EE", x"0367", x"0444", x"065B", x"0A0D", x"0CCB", x"0DD1", x"0E7A", x"0E21", x"0D37", x"0E1C", x"1038", x"1105", x"10DB", x"1090", x"0F1E", x"0D0D", x"0B84", x"096E", x"05E8", x"023F", x"FF25", x"FC5D", x"FAE0", x"FB17", x"FC33", x"FD7C", x"FE65", x"FDF1", x"FBDE", x"F8B5", x"F5C7", x"F459", x"F498", x"F58F", x"F6B2", x"F72A", x"F5E8", x"F3C1", x"F240", x"F0C1", x"EF69", x"F004", x"F206", x"F37E", x"F4E4", x"F65A", x"F60A", x"F535", x"F69A", x"F91E", x"FABB", x"FC44", x"FDB1", x"FE08", x"FFA4", x"047B", x"0A41", x"0F30", x"136B", x"15D5", x"15AD", x"1500", x"1472", x"12F8", x"1102", x"0F31", x"0CA6", x"09B7", x"07AA", x"0612", x"0476", x"038E", x"02DD", x"01AF", x"009E", x"0057", x"0042", x"010C", x"02F1", x"0511", x"06BF", x"07F8", x"07F4", x"06C2", x"05A7", x"04DC", x"046C", x"0528", x"0669", x"068A", x"05C4", x"04B3", x"0305", x"01AF", x"026B", x"03EB", x"0484", x"04E9", x"0577", x"05D7", x"0761", x"0B1B", x"0EFE", x"11C9", x"13D9", x"14CB", x"1404", x"12C2", x"119F", x"0FF1", x"0E69", x"0DA7", x"0D3B", x"0D1B", x"0DEC", x"0F4A", x"10B7", x"1281", x"1403", x"146F", x"1406", x"134F", x"1289", x"12A2", x"13FB", x"1622", x"1846", x"19C6", x"1A05", x"1982", x"1888", x"171D", x"15EE", x"15C1", x"15B5", x"15B4", x"1654", x"1681", x"157A", x"151A", x"15D9", x"15EA", x"15AF", x"1614", x"1608", x"1655", x"19B7", x"1EF3", x"2330", x"2665", x"2827", x"26F8", x"24D4", x"23F4", x"22B3", x"203C", x"1DD1", x"1AAC", x"163A", x"1319", x"1188", x"0FBA", x"0DFA", x"0CD1", x"0AA1", x"07A3", x"05AA", x"041C", x"02D9", x"0381", x"05CA", x"0839", x"0AB6", x"0C64", x"0BE9", x"0A55", x"08D1", x"075B", x"072E", x"0914", x"0AFF", x"0C43", x"0D57", x"0D27", x"0BCA", x"0C25", x"0E09", x"0F15", x"0FDA", x"10AF", x"1038", x"1015", x"12B7", x"162C", x"1843", x"19F1", x"1ABA", x"1996", x"18C9", x"195F", x"1996", x"1949", x"197C", x"193C", x"187D", x"18B2", x"19B7", x"1AAB", x"1BE6", x"1CE3", x"1C7B", x"1AD4", x"1856", x"1596", x"13C1", x"1366", x"13AF", x"146F", x"14CE", x"13B2", x"11D0", x"103B", x"0DE0", x"0B59", x"0A6F", x"0A45", x"09A3", x"0986", x"08E2", x"05C1", x"0251", x"0111", x"0079", x"FFF9", x"0096", x"0082", x"FF06", x"FF45", x"0253", x"05EA", x"0A06", x"0E89", x"1124", x"11F2", x"132F", x"1452", x"1471", x"14A1", x"146A", x"12BD", x"1101", x"1036", x"0F5D", x"0E85", x"0E11", x"0CC1", x"0A91", x"08F0", x"07BC", x"06E7", x"0770", x"08E8", x"0A04", x"0B1F", x"0BC0", x"0AB0", x"08BE", x"06CE", x"0471", x"0254", x"0222", x"02BA", x"0319", x"03D1", x"042B", x"031D", x"0255", x"02E3", x"031A", x"0292", x"0254", x"01CE", x"0130", x"0292", x"05A8", x"084B", x"0A3E", x"0BA1", x"0B71", x"0A5E", x"09EB", x"09BF", x"0955", x"0953", x"096C", x"0901", x"08E1", x"09AD", x"0ACB", x"0C5C", x"0E4B", x"0FB9", x"101C", x"0FFB", x"0F75", x"0EF7", x"0F87", x"1122", x"1319", x"14C8", x"1535", x"1416", x"1232", x"0FFB", x"0DA2", x"0BFF", x"0B4E", x"0A9D", x"0A2E", x"0A31", x"0942", x"0781", x"06C3", x"06D5", x"0679", x"0668", x"064B", x"04C3", x"0384", x"04DC", x"0773", x"0A01", x"0CF7", x"0EA6", x"0DF2", x"0CF8", x"0CE4", x"0C27", x"0AFE", x"0A22", x"0805", x"0512", x"03A5", x"0387", x"03AF", x"04F4", x"06CA", x"076D", x"0784", x"07DC", x"0737", x"0617", x"05EE", x"0624", x"063A", x"06B1", x"0641", x"040A", x"013A", x"FE78", x"FBF6", x"FB90", x"FD8F", x"0050", x"0392", x"06EA", x"0847", x"083B", x"0943", x"0A73", x"0AB0", x"0B24", x"0B09", x"08F7", x"078B", x"08CB", x"0A42", x"0B5B", x"0CED", x"0D5D", x"0BE3", x"0AED", x"0A80", x"08C7", x"06AA", x"052F", x"036F", x"0209", x"0275", x"03C1", x"053F", x"0769", x"095F", x"0A19", x"0A01", x"090E", x"074D", x"05D7", x"050B", x"0449", x"03C7", x"030A", x"013F", x"FF42", x"FD8D", x"FB4A", x"F916", x"F810", x"F72E", x"F64B", x"F682", x"F65F", x"F460", x"F2D9", x"F2C0", x"F2B6", x"F33B", x"F522", x"F5DA", x"F584", x"F728", x"FA9D", x"FDF0", x"01AA", x"053E", x"064E", x"05E8", x"05B6", x"04FC", x"0315", x"0164", x"FF45", x"FC61", x"FA20", x"F8E6", x"F812", x"F822", x"F8A7", x"F834", x"F6FC", x"F5A7", x"F3D2", x"F297", x"F30C", x"F458", x"F5BE", x"F7D2", x"F95E", x"F963", x"F8EA", x"F850", x"F6E8", x"F628", x"F70D", x"F82D", x"F917", x"FA4B", x"FA5B", x"F8D2", x"F7FC", x"F818", x"F7B4", x"F744", x"F6FB", x"F591", x"F402", x"F4C3", x"F715", x"F932", x"FB69", x"FCED", x"FC62", x"FAAF", x"F913", x"F6E8", x"F41D", x"F1F3", x"F058", x"EEFA", x"EE72", x"EEE1", x"EFEE", x"F1CF", x"F479", x"F722", x"F977", x"FB60", x"FC94", x"FDBF", x"FF97", x"0204", x"04F1", x"0836", x"0AB3", x"0B9A", x"0B4B", x"09BF", x"072C", x"04C0", x"02EE", x"010A", x"FF6A", x"FE23", x"FC2B", x"FA23", x"F992", x"FA2E", x"FB1D", x"FCB7", x"FE11", x"FDAE", x"FD4B", x"FE6C", x"001F", x"01D1", x"0408", x"0516", x"0419", x"028F", x"00BE", x"FDA8", x"FA25", x"F706", x"F38F", x"F04C", x"EE5E", x"ECFA", x"EB8C", x"EAB6", x"E999", x"E791", x"E5FF", x"E512", x"E42C", x"E421", x"E54C", x"E67F", x"E802", x"EA3E", x"EBA6", x"EB7C", x"EACA", x"E933", x"E6F9", x"E634", x"E705", x"E846", x"EA7A", x"ED1C", x"EE30", x"EEA9", x"F04B", x"F198", x"F20F", x"F2B7", x"F225", x"EF98", x"EE39", x"EF5C", x"F0CE", x"F2A5", x"F51F", x"F612", x"F57B", x"F5C6", x"F660", x"F608", x"F606", x"F647", x"F5B0", x"F539", x"F5BD", x"F620", x"F6CA", x"F838", x"F94D", x"F9BD", x"FA8C", x"FAF8", x"FABA", x"FADE", x"FAF6", x"FA38", x"F99A", x"F8F0", x"F711", x"F4D0", x"F2B3", x"F016", x"EDFA", x"ED7D", x"ED8A", x"EDD4", x"EF30", x"EFD1", x"EED8", x"EE78", x"EF10", x"EF58", x"F01B", x"F150", x"F055", x"EE31", x"EE17", x"EFC6", x"F26B", x"F6C5", x"FB57", x"FDD4", x"FF2B", x"0054", x"0042", x"FF59", x"FE99", x"FD08", x"FAA2", x"F855", x"F5A8", x"F2E0", x"F119", x"EFBE", x"EDE3", x"EC80", x"EB7A", x"EA15", x"E986", x"EA7E", x"EB73", x"ECB3", x"EF29", x"F169", x"F29E", x"F3CC", x"F42A", x"F33D", x"F2EF", x"F3EC", x"F516", x"F6E7", x"F944", x"F9AD", x"F839", x"F6EB", x"F555", x"F31F", x"F1AD", x"F01F", x"ECBD", x"E97E", x"E8AF", x"E93A", x"EB07", x"EE53", x"F14A", x"F262", x"F2EA", x"F31F", x"F25A", x"F167", x"F0FF", x"F09D", x"F06E", x"F0C6", x"F116", x"F1AB", x"F2FD", x"F467", x"F5AE", x"F753", x"F8D2", x"F99B", x"FA9D", x"FB8C", x"FB78", x"FB29", x"FB41", x"FADF", x"F9ED", x"F91D", x"F7B4", x"F5A8", x"F464", x"F3C9", x"F344", x"F348", x"F379", x"F29C", x"F1A2", x"F1C8", x"F25A", x"F350", x"F526", x"F648", x"F5DD", x"F5EE", x"F77D", x"F9B6", x"FCF2", x"00FE", x"03C4", x"04B1", x"04EF", x"041D", x"020C", x"FFC2", x"FD5E", x"FA66", x"F7A2", x"F564", x"F360", x"F25C", x"F29F", x"F2F2", x"F35D", x"F44F", x"F4C7", x"F4B2", x"F533", x"F576", x"F4AD", x"F441", x"F448", x"F388", x"F2A9", x"F21C", x"F0D0", x"EF65", x"EFAE", x"F0E1", x"F279", x"F538", x"F7B8", x"F8B0", x"F9BD", x"FB81", x"FCB9", x"FDF3", x"FF5E", x"FEB2", x"FC49", x"FAF2", x"FAC6", x"FB2F", x"FD31", x"FF6F", x"FF58", x"FDD4", x"FC21", x"F9A3", x"F74C", x"F671", x"F5C9", x"F4D5", x"F4A4", x"F486", x"F400", x"F46C", x"F569", x"F58D", x"F5D4", x"F66B", x"F5D7", x"F4A5", x"F3C2", x"F1F2", x"EF6A", x"EE34", x"EDA5", x"ECD8", x"ECC1", x"ECBB", x"EB90", x"EACB", x"EB4C", x"EBF0", x"ED41", x"EF8B", x"F0C5", x"F0E5", x"F1CF", x"F314", x"F46E", x"F727", x"FA09", x"FAC5", x"FAD2", x"FBA1", x"FC83", x"FE65", x"0216", x"0534", x"0694", x"0758", x"0727", x"05A8", x"0473", x"0395", x"01BD", x"FFD1", x"FE35", x"FBF3", x"F9F0", x"F91E", x"F813", x"F687", x"F5C7", x"F4F1", x"F3BB", x"F380", x"F3FE", x"F3D7", x"F434", x"F563", x"F617", x"F682", x"F70F", x"F645", x"F461", x"F2F4", x"F1AA", x"F092", x"F136", x"F2A8", x"F314", x"F39A", x"F467", x"F444", x"F450", x"F56C", x"F541", x"F331", x"F194", x"F0BF", x"F0AB", x"F327", x"F777", x"FAB0", x"FCB6", x"FE31", x"FE42", x"FD72", x"FD34", x"FCA6", x"FB4F", x"FA3F", x"F965", x"F843", x"F833", x"F94F", x"FA43", x"FB6F", x"FD2E", x"FE70", x"FF75", x"0149", x"0306", x"0440", x"0610", x"0806", x"095D", x"0A74", x"0B28", x"0A6E", x"092D", x"082A", x"06D2", x"05CB", x"05FF", x"0628", x"05F7", x"06BF", x"0839", x"09CE", x"0CB4", x"1050", x"11F0", x"11AE", x"1148", x"10C2", x"10EB", x"1358", x"16C9", x"18C7", x"19A0", x"1988", x"17A1", x"149C", x"1170", x"0DA3", x"093D", x"052E", x"0146", x"FDA8", x"FB42", x"F9FC", x"F96B", x"F9D4", x"FABB", x"FB3D", x"FBF9", x"FD04", x"FD7A", x"FD8E", x"FDE0", x"FDA5", x"FCCD", x"FC1F", x"FAC6", x"F866", x"F645", x"F4BA", x"F379", x"F3CF", x"F5EB", x"F7EA", x"F9E4", x"FC67", x"FE54", x"FF96", x"01C8", x"0366", x"02A0", x"00D6", x"FF64", x"FDFC", x"FE4D", x"017A", x"050D", x"077D", x"098F", x"0AD6", x"0A9E", x"0A50", x"0A37", x"0944", x"081B", x"072E", x"05E7", x"04D6", x"050B", x"05C3", x"06E6", x"08FD", x"0ADB", x"0BF8", x"0D56", x"0E66", x"0DE1", x"0CAF", x"0B46", x"08BB", x"060C", x"0442", x"0230", x"FFB0", x"FE51", x"FD67", x"FC9D", x"FCF5", x"FDCE", x"FD5F", x"FC88", x"FBE4", x"FAA3", x"F9B9", x"FA65", x"FAC1", x"F9FA", x"F98A", x"F9BC", x"FA55", x"FD2B", x"0230", x"06F8", x"0AEF", x"0E5A", x"102A", x"103E", x"0FEC", x"0EE9", x"0CF0", x"0AFA", x"0936", x"0754", x"062F", x"05DE", x"05AB", x"05B3", x"05F6", x"0596", x"04FD", x"04EE", x"04D2", x"047B", x"04A8", x"04AF", x"041C", x"037D", x"02CD", x"014D", x"FFEE", x"FF26", x"FE5C", x"FE13", x"FEC7", x"FF42", x"FF2B", x"FF55", x"FF19", x"FE1C", x"FDBE", x"FDC1", x"FC81", x"FA90", x"F917", x"F7D0", x"F7B9", x"FA6E", x"FE85", x"0200", x"04B9", x"0658", x"05D4", x"044A", x"02E7", x"012C", x"FF50", x"FE5F", x"FDF8", x"FDD3", x"FE94", x"FFEF", x"0109", x"026E", x"043E", x"05E5", x"0794", x"099E", x"0B21", x"0C0B", x"0CFC", x"0D94", x"0D80", x"0D62", x"0CE7", x"0BAD", x"0A76", x"0952", x"07B8", x"0654", x"0586", x"0441", x"02C2", x"0245", x"0261", x"0312", x"05B8", x"0913", x"0AAB", x"0AF8", x"0B3D", x"0B0F", x"0BB6", x"0F02", x"1336", x"1652", x"190E", x"1B58", x"1B8E", x"1A74", x"18F0", x"15FE", x"11FE", x"0EEF", x"0CD7", x"0B62", x"0B3D", x"0C21", x"0CF4", x"0E26", x"0FDD", x"1131", x"1210", x"1292", x"120A", x"10D7", x"0FB5", x"0E7F", x"0D67", x"0CFE", x"0CB9", x"0C4E", x"0C36", x"0BDF", x"0AF1", x"0ACE", x"0B6E", x"0B9D", x"0C2B", x"0D88", x"0E74", x"0F89", x"11FB", x"138D", x"1280", x"108B", x"0E6F", x"0BCE", x"0AE9", x"0C9A", x"0E35", x"0EDA", x"0FD2", x"103C", x"0FA1", x"0F83", x"0FD4", x"0F72", x"0F23", x"0F58", x"0F33", x"0F48", x"1008", x"1091", x"1107", x"11EE", x"1258", x"127C", x"134F", x"13E3", x"1360", x"12A9", x"114F", x"0E87", x"0C1B", x"0AB1", x"0913", x"07C5", x"0795", x"06DF", x"05DB", x"0617", x"0640", x"04FC", x"0403", x"039D", x"0324", x"0491", x"089F", x"0C08", x"0DCD", x"0F3A", x"0FC7", x"0F88", x"112C", x"148A", x"1780", x"1A65", x"1DC8", x"1FF5", x"20DB", x"213C", x"2056", x"1DD0", x"1AE5", x"17BD", x"1429", x"1114", x"0E93", x"0C24", x"0A75", x"0995", x"08FD", x"0915", x"0A2C", x"0B1D", x"0BB1", x"0C51", x"0C58", x"0B93", x"0B02", x"0A7D", x"0972", x"08A3", x"07FD", x"070B", x"0655", x"069F", x"06F0", x"0792", x"08F3", x"0A44", x"0B2F", x"0C4D", x"0CDD", x"0B78", x"08D9", x"05F1", x"02F1", x"0155", x"0276", x"053D", x"085F", x"0B87", x"0DA8", x"0DC4", x"0C7F", x"0A82", x"07CC", x"053E", x"03BE", x"0335", x"0398", x"0552", x"0784", x"09C0", x"0C35", x"0EDA", x"116A", x"1474", x"17F3", x"1B03", x"1D77", x"1F55", x"1FF3", x"1F88", x"1EB6", x"1D8A", x"1BF8", x"1ABA", x"1995", x"180E", x"16E4", x"1619", x"14CB", x"139D", x"1341", x"133B", x"13E3", x"162D", x"1872", x"18B6", x"17A1", x"15B9", x"12E4", x"1122", x"1214", x"13DD", x"153F", x"1708", x"1821", x"1745", x"1581", x"130D", x"0E63", x"08C1", x"0436", x"009D", x"FE08", x"FDA1", x"FE7C", x"FF32", x"00CE", x"035D", x"0564", x"06C0", x"0796", x"06D9", x"04DE", x"02FA", x"014A", x"FFBA", x"FEFC", x"FEC1", x"FE9A", x"FEC9", x"FED2", x"FE80", x"FE8B", x"FF24", x"FFC4", x"0122", x"0386", x"05AF", x"0811", x"0B04", x"0C64", x"0B16", x"088B", x"052E", x"0189", x"003C", x"0226", x"050B", x"0889", x"0CA0", x"0F96", x"10A3", x"110A", x"1032", x"0DC4", x"0B61", x"09E5", x"08C2", x"08B0", x"09C8", x"0ABD", x"0B8B", x"0C9A", x"0D27", x"0D3D", x"0D63", x"0CFD", x"0B94", x"09D1", x"0724", x"0376", x"004D", x"FDFB", x"FC1A", x"FB9E", x"FC37", x"FC2F", x"FC23", x"FCEF", x"FCC9", x"FB50", x"FA0B", x"F840", x"F5DA", x"F58F", x"F790", x"F908", x"FA03", x"FB35", x"FB57", x"FB5B", x"FDE5", x"01F1", x"057C", x"094B", x"0CC1", x"0E18", x"0E09", x"0D44", x"0A84", x"066F", x"02D9", x"FFBA", x"FD2C", x"FC46", x"FC50", x"FC30", x"FC94", x"FDA5", x"FE94", x"FFEF", x"01F8", x"0390", x"04BE", x"05FB", x"06DC", x"076E", x"0887", x"09D3", x"0B11", x"0CA3", x"0DDB", x"0DE5", x"0D58", x"0C36", x"0A1B", x"07F4", x"0687", x"0528", x"0433", x"0444", x"0413", x"0270", x"FFF6", x"FCAA", x"F8E3", x"F689", x"F6A6", x"F844", x"FABE", x"FD7A", x"FEDC", x"FE7D", x"FCF9", x"FA78", x"F769", x"F4FE", x"F391", x"F2D2", x"F31F", x"F43F", x"F545", x"F640", x"F754", x"F80A", x"F89F", x"F9CA", x"FB22", x"FC93", x"FE40", x"FF6A", x"FFA5", x"FF32", x"FE0F", x"FC00", x"FA0A", x"F838", x"F5E4", x"F384", x"F1C1", x"EFED", x"EE42", x"EDD9", x"EE19", x"EE6E", x"F049", x"F3B3", x"F6E0", x"F940", x"FAB6", x"FA06", x"F7EC", x"F71A", x"F82E", x"FA51", x"FD76", x"0107", x"031B", x"0398", x"0336", x"0170", x"FE07", x"FA85", x"F79C", x"F53F", x"F40F", x"F42F", x"F4C9", x"F569", x"F6A3", x"F84C", x"F9C0", x"FAD6", x"FB50", x"FAB8", x"F921", x"F725", x"F543", x"F37F", x"F1FE", x"F13D", x"F145", x"F183", x"F1B7", x"F1F2", x"F1E0", x"F19A", x"F200", x"F365", x"F524", x"F703", x"F96C", x"FB84", x"FC75", x"FC15", x"FA4E", x"F6F0", x"F369", x"F181", x"F1BD", x"F38D", x"F695", x"FA0B", x"FC99", x"FDDE", x"FE17", x"FD32", x"FB77", x"F9BB", x"F8B6", x"F825", x"F7A4", x"F74D", x"F702", x"F69B", x"F634", x"F610", x"F5BE", x"F4DF", x"F3FB", x"F362", x"F289", x"F133", x"EFAD", x"EDB8", x"EB67", x"EA17", x"EA53", x"EB2F", x"EC4C", x"EDB0", x"EE60", x"EDE3", x"ED35", x"ECA4", x"EBBA", x"EB7A", x"ECFD", x"EF5F", x"F174", x"F2F8", x"F31B", x"F14E", x"EF74", x"EF47", x"F0D1", x"F3AB", x"F7DB", x"FC21", x"FF16", x"00AE", x"00D8", x"FF0F", x"FBDE", x"F875", x"F519", x"F1CD", x"EEE6", x"EC6D", x"EA53", x"E90D", x"E8DB", x"E989", x"EA8C", x"EBA7", x"EC64", x"ECB7", x"ECA6", x"EC4D", x"EBD2", x"EB42", x"EADC", x"EAC8", x"EB41", x"EBFB", x"ECCE", x"ED5F", x"ED67", x"ECC7", x"EC1B", x"EB90", x"EB67", x"EBE7", x"ECF9", x"EDC6", x"ED91", x"EC5A", x"EA19", x"E7A8", x"E693", x"E7B8", x"EAF8", x"EF6F", x"F44E", x"F800", x"F9A3", x"F90D", x"F6B5", x"F358", x"F003", x"EDB1", x"ECBF", x"ECD0", x"ED72", x"EE90", x"F015", x"F1E9", x"F450", x"F758", x"FA6F", x"FD36", x"FFA9", x"014E", x"01B2", x"0138", x"FFF2", x"FDF5", x"FC01", x"FB06", x"FAA6", x"FAA0", x"FB25", x"FB2B", x"FA1D", x"F8C8", x"F7A9", x"F641", x"F573", x"F66C", x"F885", x"FB1C", x"FE2D", x"006A", x"0066", x"FF3E", x"FEB0", x"FEE4", x"0031", x"02B0", x"04E8", x"0557", x"041F", x"017F", x"FD6F", x"F8AA", x"F420", x"F03B", x"ED20", x"EB2D", x"EA3F", x"EA41", x"EAFA", x"EC54", x"EE0E", x"EFAE", x"F0AB", x"F0D5", x"F039", x"EEE4", x"ED2E", x"EBC1", x"EA5F", x"E92F", x"E8C4", x"E90C", x"E99A", x"EA8B", x"EBB2", x"EC36", x"EC80", x"ED8A", x"EF1D", x"F0F9", x"F3A3", x"F6DB", x"F984", x"FB59", x"FC17", x"FAF1", x"F81C", x"F54C", x"F3E1", x"F48E", x"F6FF", x"FA98", x"FE05", x"FFFF", x"FFDA", x"FE2C", x"FB9F", x"F8AC", x"F65F", x"F5C9", x"F5FB", x"F5D0", x"F5CB", x"F601", x"F5BF", x"F5AA", x"F642", x"F61B", x"F4C1", x"F38D", x"F2BF", x"F1A4", x"F0F2", x"F06B", x"EEA0", x"EC17", x"EA50", x"E944", x"E8CE", x"E9AA", x"EAD2", x"EAC6", x"EA1A", x"E955", x"E7CE", x"E623", x"E5A1", x"E61E", x"E71E", x"E8EC", x"EABF", x"EB3F", x"EA9F", x"EA26", x"EAC0", x"ECEF", x"F0E6", x"F60F", x"FB1E", x"FED8", x"00A2", x"00A7", x"FF06", x"FC55", x"F9E6", x"F85A", x"F728", x"F61F", x"F59B", x"F58A", x"F59F", x"F66F", x"F7B8", x"F8A7", x"F901", x"F937", x"F949", x"F942", x"F993", x"FA3B", x"FB14", x"FC13", x"FD05", x"FDC5", x"FE59", x"FE85", x"FE06", x"FCCF", x"FAE4", x"F87E", x"F670", x"F57A", x"F5AA", x"F6AB", x"F7BD", x"F7B7", x"F635", x"F369", x"F00A", x"ED6C", x"ECDC", x"EE64", x"F161", x"F55D", x"F906", x"FAD1", x"FA9F", x"F8E6", x"F5BB", x"F21D", x"EFB9", x"EEAE", x"EE19", x"EDF1", x"EE4C", x"EE67", x"EEA1", x"EFC8", x"F18E", x"F361", x"F597", x"F84A", x"FACC", x"FCEF", x"FEB3", x"FF70", x"FEFB", x"FE02", x"FCC9", x"FB97", x"FB01", x"FB1C", x"FB1B", x"FAAA", x"FA11", x"F8F5", x"F796", x"F725", x"F810", x"F9CF", x"FC6A", x"FF81", x"0183", x"019A", x"0105", x"00B8", x"015F", x"03DF", x"0817", x"0BF3", x"0E23", x"0EB3", x"0DC5", x"0B7E", x"08F3", x"06B7", x"0488", x"0293", x"0128", x"0020", x"FF7C", x"FFA7", x"0074", x"01B0", x"032A", x"045F", x"04BD", x"044D", x"030B", x"0102", x"FE9A", x"FC41", x"FA07", x"F822", x"F6D0", x"F615", x"F5FB", x"F690", x"F751", x"F803", x"F89D", x"F8FE", x"F92F", x"F9CC", x"FAED", x"FC01", x"FCDC", x"FD1A", x"FBD6", x"F925", x"F67B", x"F516", x"F595", x"F84F", x"FCAC", x"00F0", x"03CE", x"0520", x"050F", x"03FD", x"029A", x"0213", x"02B2", x"03EE", x"0568", x"0719", x"088B", x"0974", x"0A77", x"0B87", x"0B8D", x"0AB4", x"09F1", x"094E", x"08A2", x"087A", x"083D", x"0695", x"042C", x"0212", x"0019", x"FE9B", x"FE71", x"FEB6", x"FE61", x"FE35", x"FE4C", x"FDC7", x"FD2C", x"FD91", x"FE3C", x"FF03", x"00AA", x"0232", x"020C", x"00E0", x"FFD8", x"FF5F", x"005B", x"0394", x"07CE", x"0B4A", x"0DA1", x"0E73", x"0D66", x"0AF8", x"081B", x"0542", x"02CD", x"00ED", x"FF52", x"FDFB", x"FCCE", x"FBD3", x"FAFA", x"FA6A", x"F98A", x"F846", x"F714", x"F5F0", x"F49F", x"F35C", x"F280", x"F1BB", x"F14F", x"F191", x"F25F", x"F364", x"F4D5", x"F672", x"F78C", x"F7F0", x"F7C9", x"F72D", x"F6C0", x"F750", x"F8DE", x"FAC4", x"FC83", x"FD32", x"FC3D", x"FA1E", x"F855", x"F7D8", x"F93A", x"FC91", x"011E", x"0541", x"0812", x"093D", x"08B6", x"06CC", x"04C7", x"03D0", x"03E5", x"049B", x"05E5", x"078D", x"095B", x"0B94", x"0EB8", x"120D", x"14C4", x"1719", x"1920", x"1A4C", x"1ABA", x"1ABF", x"1A33", x"18E8", x"17B2", x"16B5", x"159F", x"14D6", x"1488", x"140D", x"1320", x"11F9", x"1049", x"0E0D", x"0C99", x"0C2F", x"0C96", x"0E11", x"104C", x"114B", x"108D", x"0F04", x"0D35", x"0BDF", x"0C8D", x"0EC2", x"1070", x"10CC", x"0FF6", x"0D6C", x"09B4", x"064C", x"034D", x"008A", x"FE67", x"FCC8", x"FB2A", x"F9F5", x"F9AD", x"F9EB", x"FAB7", x"FC11", x"FD04", x"FD5C", x"FD6D", x"FCCC", x"FB42", x"F99D", x"F81B", x"F681", x"F52B", x"F483", x"F414", x"F42F", x"F55A", x"F6F8", x"F8A1", x"FA42", x"FB8B", x"FC7D", x"FDC3", x"FF72", x"0138", x"0342", x"0527", x"05C6", x"0541", x"048F", x"040A", x"046F", x"069C", x"09D1", x"0C92", x"0E9D", x"0FD5", x"0FE4", x"0EEF", x"0DCD", x"0CB6", x"0BDA", x"0B71", x"0B81", x"0BC2", x"0C22", x"0C87", x"0D28", x"0DBA", x"0DA2", x"0CC7", x"0BE2", x"0AD6", x"09BC", x"090E", x"087B", x"0735", x"058F", x"0419", x"024A", x"0089", x"FFA6", x"FF13", x"FE51", x"FE0A", x"FDCD", x"FCD2", x"FBC4", x"FB64", x"FB11", x"FB75", x"FD54", x"FF53", x"0004", x"FFF7", x"FF83", x"FEAB", x"FF0D", x"018F", x"04CA", x"07AA", x"0A3F", x"0BB8", x"0B6D", x"09F2", x"07F5", x"0598", x"039F", x"02B8", x"028E", x"02D2", x"035F", x"03FA", x"04BC", x"05B7", x"06AF", x"0790", x"08D7", x"0A27", x"0B6C", x"0CED", x"0EA2", x"0FF5", x"1136", x"127C", x"1333", x"1376", x"13EB", x"144B", x"1460", x"1447", x"13A2", x"11CD", x"0F7C", x"0D91", x"0C3F", x"0BD1", x"0C5F", x"0C6A", x"0AA0", x"0786", x"03E8", x"00B2", x"FF12", x"FFD6", x"01E4", x"0405", x"05D4", x"06C2", x"061A", x"0465", x"028B", x"013C", x"007D", x"0086", x"0109", x"018C", x"0201", x"02F5", x"04BD", x"06F5", x"0946", x"0BD2", x"0E4F", x"1040", x"1198", x"127D", x"126C", x"1173", x"1034", x"0EE7", x"0D58", x"0C2F", x"0BC8", x"0B91", x"0B7F", x"0B99", x"0B06", x"097D", x"07F2", x"06E6", x"0671", x"0755", x"095D", x"0AB8", x"0ADB", x"0A8E", x"0A24", x"0A38", x"0C02", x"0F1F", x"11ED", x"13D8", x"1500", x"14B4", x"1334", x"117E", x"0FC5", x"0E34", x"0D33", x"0C93", x"0BF7", x"0B97", x"0B91", x"0B95", x"0C05", x"0C9B", x"0CB7", x"0C8A", x"0C72", x"0B9A", x"09E6", x"081B", x"0614", x"03B5", x"01D8", x"00B2", x"FFAF", x"FF64", x"006C", x"0211", x"0403", x"0643", x"07D0", x"084B", x"086C", x"087B", x"0839", x"087F", x"08F5", x"085A", x"06CB", x"054D", x"03F5", x"0367", x"04B2", x"071B", x"095C", x"0B6F", x"0D39", x"0DD8", x"0D7A", x"0CC2", x"0BD2", x"0B16", x"0B1F", x"0BBB", x"0C74", x"0D38", x"0D8E", x"0D7E", x"0D4E", x"0CE9", x"0C40", x"0C10", x"0C46", x"0C49", x"0C5A", x"0CA8", x"0CA1", x"0C51", x"0C0E", x"0B3C", x"09E7", x"08F4", x"08A0", x"08EC", x"0A4A", x"0C1A", x"0D36", x"0DB4", x"0DB4", x"0CE1", x"0C3C", x"0CE2", x"0D91", x"0D4F", x"0C6F", x"0ACC", x"0863", x"072E", x"080F", x"09A3", x"0B42", x"0D0F", x"0DD4", x"0CFF", x"0B7E", x"0969", x"06BC", x"048D", x"037B", x"02FF", x"030E", x"03A1", x"03F7", x"041C", x"04A7", x"0521", x"056E", x"05FF", x"0652", x"05B6", x"04DF", x"0424", x"0335", x"028D", x"0268", x"0213", x"0199", x"01A8", x"0207", x"028D", x"0356", x"03A5", x"02B9", x"0141", x"FFC9", x"FE6D", x"FE67", x"000C", x"0174", x"0192", x"00BC", x"FEE4", x"FCBC", x"FC67", x"FE4C", x"00C8", x"0342", x"05A4", x"06DD", x"068E", x"05C7", x"04B3", x"0367", x"02C4", x"0323", x"040E", x"0540", x"06CC", x"088D", x"0A99", x"0CD6", x"0ECA", x"1072", x"11DC", x"12A7", x"1309", x"133A", x"12C6", x"1194", x"1055", x"0ED8", x"0CEA", x"0B5A", x"0A4D", x"0958", x"091D", x"09EC", x"0A78", x"0A82", x"0ABE", x"0AB8", x"0A99", x"0C2C", x"0F1E", x"1157", x"12AB", x"138F", x"1325", x"1259", x"1317", x"1459", x"1474", x"140D", x"1340", x"111F", x"0E75", x"0C1E", x"0965", x"065C", x"041A", x"0263", x"00AB", x"FF73", x"FE59", x"FD12", x"FC35", x"FBE1", x"FB6E", x"FB72", x"FBDD", x"FB93", x"FAAF", x"F9BA", x"F810", x"F60F", x"F4E6", x"F415", x"F327", x"F305", x"F3DF", x"F503", x"F73B", x"FA7C", x"FD15", x"FEBD", x"0032", x"00DE", x"0145", x"02F5", x"0551", x"068E", x"0735", x"0747", x"0637", x"0536", x"05B6", x"06A6", x"0760", x"0863", x"08EA", x"07F1", x"0615", x"0371", x"000D", x"FCF9", x"FAD7", x"F966", x"F8E0", x"F92E", x"F95C", x"F9AD", x"FA41", x"FA21", x"F990", x"F9C6", x"FA10", x"FA02", x"FA83", x"FB3C", x"FB26", x"FB36", x"FBAC", x"FAEF", x"F924", x"F780", x"F594", x"F40D", x"F481", x"F601", x"F6DA", x"F753", x"F724", x"F569", x"F43F", x"F4F6", x"F5FD", x"F68D", x"F723", x"F68E", x"F4F7", x"F506", x"F71F", x"F99D", x"FC9B", x"FFA8", x"00F3", x"00BE", x"004E", x"FF0D", x"FD2C", x"FC29", x"FBBF", x"FB74", x"FC2E", x"FD7F", x"FE15", x"FE82", x"FF0C", x"FECF", x"FE6D", x"FEF6", x"FF67", x"FF45", x"FF72", x"FFAF", x"FF4C", x"FF1A", x"FF05", x"FE2E", x"FD13", x"FC69", x"FBCC", x"FB5E", x"FB31", x"FA34", x"F846", x"F609", x"F341", x"F082", x"EF5E", x"EF99", x"EFCE", x"EFF3", x"EF5A", x"ECF8", x"EA65", x"E9C7", x"EAC3", x"ECC1", x"EFCA", x"F24F", x"F2D4", x"F233", x"F0DC", x"EE56", x"EBA5", x"E9A8", x"E7F0", x"E6B5", x"E6F2", x"E7C5", x"E8FD", x"EAF3", x"ECEE", x"EE19", x"EF42", x"F088", x"F131", x"F1C2", x"F2A5", x"F2EE", x"F2D9", x"F331", x"F34E", x"F2FF", x"F332", x"F35C", x"F327", x"F3B9", x"F4F8", x"F5D0", x"F6C3", x"F7DB", x"F77A", x"F684", x"F6FB", x"F7DA", x"F82A", x"F8F0", x"F968", x"F85B", x"F836", x"FA9F", x"FD85", x"001D", x"0319", x"04EA", x"0483", x"03CB", x"02D7", x"0079", x"FDE2", x"FC9B", x"FBEB", x"FBC7", x"FCA9", x"FD3C", x"FCBE", x"FC23", x"FB65", x"FA4A", x"F977", x"F8AF", x"F722", x"F538", x"F360", x"F123", x"EF36", x"EE17", x"ECFC", x"EC21", x"EC08", x"EC2A", x"EC7A", x"EDD1", x"EF68", x"F037", x"F0F5", x"F123", x"EFD2", x"EEAB", x"EEE4", x"EF11", x"EF04", x"EF46", x"EE67", x"EC35", x"EB6D", x"EC76", x"EDF7", x"F04B", x"F342", x"F4DB", x"F534", x"F596", x"F542", x"F458", x"F432", x"F4BD", x"F55F", x"F70B", x"F947", x"FB0F", x"FD1A", x"FF11", x"FF93", x"FF6C", x"FF6C", x"FE62", x"FCF7", x"FC67", x"FBAB", x"FA64", x"FA67", x"FB05", x"FA5B", x"F963", x"F84C", x"F5F1", x"F3FC", x"F46A", x"F57B", x"F65F", x"F7CE", x"F83D", x"F6FC", x"F6AB", x"F7B8", x"F81B", x"F833", x"F806", x"F5D5", x"F307", x"F2B6", x"F43D", x"F6A1", x"FA60", x"FDEA", x"FF46", x"FFAE", x"FFF0", x"FEB8", x"FD1A", x"FBF6", x"FA7C", x"F8FF", x"F8C0", x"F8CA", x"F851", x"F825", x"F76C", x"F53E", x"F30B", x"F131", x"EEC3", x"EC66", x"EAD3", x"E8AF", x"E665", x"E4FB", x"E3B5", x"E22A", x"E153", x"E0FF", x"E083", x"E0F7", x"E202", x"E2B5", x"E39E", x"E4D6", x"E558", x"E5EA", x"E791", x"E93A", x"EAC0", x"ECC6", x"ED9B", x"EC97", x"EBD1", x"EC3D", x"ED1E", x"EF99", x"F32F", x"F54B", x"F59C", x"F5B6", x"F4DC", x"F320", x"F242", x"F1B9", x"F097", x"F077", x"F20C", x"F40C", x"F6C0", x"FA69", x"FD2C", x"FEBD", x"0062", x"0197", x"01CC", x"01FE", x"0225", x"0164", x"00B8", x"009B", x"001B", x"FF9B", x"FF75", x"FEF8", x"FE5A", x"FE86", x"FECB", x"FEF3", x"FFDC", x"0083", x"FFFC", x"FFBE", x"003B", x"0082", x"0145", x"02CD", x"02E2", x"016E", x"00D8", x"0129", x"0191", x"0322", x"04F9", x"04B5", x"02CB", x"00D3", x"FDDF", x"F9EE", x"F6BD", x"F43F", x"F1D9", x"F0D1", x"F136", x"F157", x"F100", x"F0CB", x"F02B", x"EF32", x"EEAF", x"EE14", x"ECD9", x"EB6E", x"EA1B", x"E8D6", x"E7E5", x"E728", x"E643", x"E58B", x"E529", x"E4FA", x"E5B0", x"E731", x"E8D8", x"EAE9", x"ED9E", x"EFB1", x"F0FB", x"F2C7", x"F4D2", x"F656", x"F839", x"F9E1", x"F97B", x"F83B", x"F86E", x"F9BA", x"FBD6", x"FF51", x"0267", x"030E", x"0269", x"0177", x"FF70", x"FD14", x"FB9E", x"FA6B", x"F95D", x"F9A1", x"FAC6", x"FBC4", x"FD10", x"FE53", x"FEBF", x"FEC9", x"FECC", x"FE3C", x"FDA3", x"FDA7", x"FD96", x"FD88", x"FDE7", x"FDD8", x"FCE2", x"FBF0", x"FAA3", x"F8B4", x"F77D", x"F742", x"F6FD", x"F71C", x"F7C1", x"F736", x"F5E6", x"F58B", x"F58D", x"F54C", x"F5B5", x"F5DC", x"F448", x"F315", x"F428", x"F665", x"F9DB", x"FEB3", x"026A", x"03C0", x"045D", x"0459", x"02D3", x"014B", x"0055", x"FF0D", x"FE47", x"FF4F", x"00C4", x"022A", x"03F7", x"051B", x"04EB", x"04E0", x"0514", x"04DE", x"0524", x"060E", x"067F", x"06E4", x"0817", x"0912", x"09B6", x"0AB0", x"0B4C", x"0AFE", x"0AB7", x"0A34", x"08EE", x"07B1", x"06C7", x"0556", x"0434", x"03C7", x"02EF", x"01CC", x"00B0", x"FE8E", x"FB5B", x"F956", x"F8BF", x"F94F", x"FBC6", x"FF29", x"00EC", x"011D", x"00BA", x"FEE1", x"FC25", x"FA30", x"F875", x"F67C", x"F600", x"F6FF", x"F83E", x"FA0F", x"FC84", x"FE09", x"FEDA", x"0013", x"00F6", x"013A", x"01CE", x"027A", x"02A5", x"0351", x"0458", x"04D5", x"0500", x"04F8", x"045D", x"03B4", x"03AA", x"0393", x"03B5", x"046E", x"0499", x"0400", x"03AA", x"0337", x"0266", x"0299", x"0354", x"02B9", x"01C1", x"020E", x"02EC", x"04F5", x"0948", x"0D74", x"0F2D", x"0FBD", x"0FAA", x"0E01", x"0C32", x"0B96", x"0A99", x"0950", x"09AC", x"0AEE", x"0B85", x"0C2E", x"0CA2", x"0BAE", x"0A4E", x"09BE", x"08F3", x"078C", x"0656", x"0505", x"037B", x"0281", x"0212", x"0179", x"00F3", x"0090", x"004A", x"006A", x"00E2", x"012B", x"01A2", x"0246", x"025F", x"025D", x"02E2", x"0323", x"02FF", x"0334", x"0296", x"0059", x"FE2D", x"FD88", x"FE0B", x"0066", x"049A", x"0816", x"098C", x"0A36", x"0A42", x"094B", x"088C", x"088E", x"085E", x"0870", x"09D5", x"0BC9", x"0D77", x"0F30", x"107F", x"10B7", x"105E", x"0FAA", x"0E89", x"0D59", x"0CC6", x"0CBA", x"0D2E", x"0D9D", x"0D7C", x"0CF9", x"0C4E", x"0B78", x"0AEC", x"0AFE", x"0AEE", x"0AE0", x"0BA3", x"0C5F", x"0C32", x"0BC3", x"0B2B", x"097B", x"07AF", x"0684", x"046B", x"0130", x"FF07", x"FE52", x"FEDE", x"01B5", x"0614", x"0909", x"0A42", x"0AD4", x"0A24", x"086C", x"0759", x"06CB", x"05E9", x"0618", x"07AB", x"0914", x"0A23", x"0AEB", x"0A5F", x"0886", x"070C", x"05FC", x"04A5", x"03DA", x"0355", x"0237", x"00F8", x"005B", x"FF7A", x"FE49", x"FD65", x"FC77", x"FB57", x"FAD3", x"FACA", x"FAB9", x"FB06", x"FBB7", x"FC61", x"FD67", x"FF04", x"0062", x"0152", x"0202", x"01BD", x"00CF", x"00D9", x"0236", x"04BA", x"0893", x"0CE6", x"0FE0", x"1156", x"11C3", x"10C4", x"0ED9", x"0D5C", x"0C68", x"0BF7", x"0CF3", x"0EF5", x"10DF", x"129B", x"140F", x"147F", x"1444", x"1416", x"1385", x"1254", x"1141", x"1055", x"0F71", x"0F31", x"0F70", x"0F70", x"0EF8", x"0E58", x"0DA3", x"0D63", x"0DB1", x"0E64", x"0F8E", x"1106", x"1214", x"12F3", x"13EB", x"1444", x"1459", x"1522", x"1596", x"1481", x"1353", x"12D6", x"12CE", x"14A0", x"18C9", x"1C1A", x"1CC1", x"1BD9", x"1919", x"1442", x"0FFE", x"0D0C", x"09D0", x"074C", x"0757", x"084B", x"0921", x"0AA4", x"0B43", x"0974", x"074D", x"0638", x"04CB", x"037D", x"0331", x"02A0", x"0164", x"0149", x"01DC", x"01C0", x"018E", x"01D0", x"021B", x"02FE", x"050B", x"0772", x"09CA", x"0C3B", x"0E88", x"10C4", x"1328", x"1509", x"1640", x"16F9", x"165B", x"1418", x"11E5", x"109B", x"1077", x"124E", x"15AD", x"17E7", x"1818", x"1703", x"1485", x"10D9", x"0DB9", x"0B66", x"094F", x"0846", x"08B9", x"0981", x"09F7", x"0A3F", x"09CA", x"087D", x"071C", x"05EA", x"04C4", x"0405", x"03F0", x"049B", x"05B0", x"06A9", x"0731", x"077D", x"074F", x"06FA", x"0721", x"071F", x"0606", x"0509", x"04C7", x"045E", x"0411", x"04AB", x"0496", x"0362", x"0306", x"034B", x"0208", x"0026", x"FF0C", x"FE15", x"FE7D", x"0263", x"07C5", x"0BB6", x"0E72", x"0FEE", x"0EF3", x"0CF6", x"0BEF", x"0B04", x"0A55", x"0BAF", x"0E86", x"1132", x"13BB", x"15C0", x"15DA", x"14DC", x"1456", x"13F1", x"1347", x"130F", x"12E9", x"121E", x"1180", x"1166", x"10EF", x"0FD4", x"0E6D", x"0CB3", x"0A9B", x"08C7", x"075A", x"05F9", x"04C8", x"0405", x"03B9", x"03DE", x"043A", x"0469", x"040A", x"02EE", x"00F3", x"FEB0", x"FD26", x"FCF8", x"FE62", x"011E", x"044A", x"0656", x"06A6", x"0530", x"021F", x"FDFF", x"FA11", x"F75A", x"F619", x"F63F", x"F77A", x"F8C7", x"F989", x"F9F3", x"FA5D", x"FADD", x"FB92", x"FC87", x"FD72", x"FE4A", x"FF89", x"0136", x"0309", x"04E0", x"0659", x"0704", x"0734", x"07A5", x"087A", x"0957", x"0A75", x"0BA9", x"0C52", x"0C95", x"0D1B", x"0D9A", x"0DAE", x"0E38", x"0F5C", x"0FC1", x"0EF1", x"0DE5", x"0CA2", x"0BAA", x"0CE3", x"1035", x"1313", x"1469", x"148B", x"129B", x"0EE8", x"0BB9", x"0963", x"06E8", x"05B6", x"06C4", x"086B", x"0A0D", x"0BEF", x"0C60", x"0A52", x"081F", x"069F", x"04C0", x"0331", x"0292", x"0155", x"FF7C", x"FEF4", x"FEFB", x"FE08", x"FCD8", x"FBF7", x"FAA3", x"F9A9", x"F9FD", x"FA8D", x"FA7F", x"FA8E", x"FAFC", x"FB7A", x"FC21", x"FCCF", x"FCE3", x"FC28", x"FA5A", x"F7A7", x"F514", x"F363", x"F372", x"F630", x"FADB", x"FF61", x"0297", x"0470", x"0410", x"0231", x"006B", x"FF4A", x"FEC1", x"FFFE", x"0309", x"0665", x"095E", x"0BC4", x"0CDB", x"0CC5", x"0CCF", x"0D26", x"0D9D", x"0E52", x"0F5F", x"1046", x"10EB", x"1126", x"10CC", x"0FAB", x"0E0F", x"0C97", x"0BC8", x"0B01", x"09D0", x"08CE", x"07A0", x"05D3", x"0417", x"02BF", x"003C", x"FD2C", x"FB65", x"F9FE", x"F797", x"F564", x"F3BB", x"F1EE", x"F234", x"F680", x"FC23", x"009B", x"0439", x"05BE", x"03E0", x"00E0", x"FE56", x"FB4F", x"F8B1", x"F88B", x"F9BE", x"FAB2", x"FB9B", x"FB7F", x"F91E", x"F5D5", x"F302", x"F049", x"ED8A", x"EB73", x"E968", x"E742", x"E5EC", x"E577", x"E543", x"E53A", x"E53C", x"E520", x"E4EE", x"E4AA", x"E422", x"E372", x"E2AA", x"E1F5", x"E213", x"E329", x"E49F", x"E6B3", x"E95C", x"EB62", x"EC26", x"EC74", x"ECB1", x"ED76", x"F067", x"F5AF", x"FB72", x"0015", x"0316", x"0379", x"014D", x"FDEC", x"FAAA", x"F813", x"F72E", x"F839", x"FA69", x"FC8D", x"FDEE", x"FE43", x"FDEA", x"FD1C", x"FC34", x"FB8B", x"FB1B", x"FAD1", x"FB0B", x"FC12", x"FCFF", x"FDD1", x"FEAE", x"FF2D", x"FF24", x"FF7F", x"0009", x"001D", x"0035", x"00D3", x"00CF", x"0088", x"00BC", x"00B3", x"0025", x"0092", x"01B4", x"01C6", x"00D0", x"FF54", x"FC9E", x"FA1F", x"FA46", x"FC81", x"FEB1", x"0083", x"00EB", x"FE8E", x"FA7E", x"F6A3", x"F2D8", x"EF8D", x"EE2C", x"EE44", x"EEC7", x"EF9A", x"F01F", x"EF12", x"ECEA", x"EAAD", x"E865", x"E67D", x"E59B", x"E50E", x"E449", x"E3A7", x"E323", x"E28E", x"E250", x"E2A0", x"E327", x"E417", x"E57F", x"E6FC", x"E86E", x"E9C1", x"EAB0", x"EB9F", x"ECF5", x"EE70", x"EFFD", x"F1F9", x"F368", x"F357", x"F219", x"EFDB", x"ECF2", x"EB3F", x"EC60", x"EF6D", x"F339", x"F6EB", x"F8EA", x"F843", x"F62B", x"F3B7", x"F162", x"F01C", x"F091", x"F1FE", x"F388", x"F4AA", x"F4A0", x"F33C", x"F10D", x"EE91", x"EC4B", x"EAC6", x"E9F4", x"E9B9", x"EA1D", x"EA99", x"EA9A", x"EA79", x"EA1C", x"E950", x"E8F5", x"E963", x"E9C4", x"EA30", x"EB34", x"EBF0", x"EC2B", x"ED01", x"EDD5", x"ED8E", x"ED84", x"EE53", x"EE77", x"EDC8", x"ED04", x"EB12", x"E859", x"E80A", x"EB0F", x"EF99", x"F528", x"FAA3", x"FD56", x"FD2F", x"FC4B", x"FB0D", x"F98B", x"F989", x"FB34", x"FD36", x"FF56", x"013D", x"018D", x"0031", x"FE8A", x"FCD8", x"FB95", x"FB82", x"FC10", x"FC82", x"FCEC", x"FD1F", x"FCCE", x"FC92", x"FC91", x"FC6C", x"FC73", x"FCE4", x"FCFD", x"FCDE", x"FCF9", x"FCA8", x"FBE6", x"FBA8", x"FB90", x"FB34", x"FBA0", x"FCC5", x"FCE0", x"FBD5", x"F9CD", x"F64E", x"F29C", x"F17F", x"F327", x"F615", x"F97D", x"FBD0", x"FB13", x"F7A1", x"F336", x"EE4E", x"E9F2", x"E78F", x"E73D", x"E82A", x"EA12", x"EC29", x"EDDF", x"EF57", x"F0B0", x"F1E5", x"F33E", x"F4AB", x"F5BB", x"F6E7", x"F81E", x"F892", x"F8B3", x"F92B", x"F983", x"F9FB", x"FB9B", x"FD74", x"FEA0", x"001A", x"01A7", x"021C", x"0246", x"02B9", x"021B", x"010F", x"01A3", x"02F9", x"03B3", x"0473", x"041D", x"016C", x"FECB", x"FEAF", x"000E", x"024E", x"0521", x"05F0", x"0351", x"FF6D", x"FB54", x"F725", x"F4A2", x"F4A1", x"F5B4", x"F79F", x"FA7F", x"FCB7", x"FDB1", x"FE38", x"FDCC", x"FC5B", x"FB56", x"FAC0", x"F9F3", x"F964", x"F8E8", x"F718", x"F4C1", x"F2E6", x"F0FF", x"EF7E", x"EF49", x"EF5E", x"EEED", x"EEE7", x"EEB4", x"ED84", x"EC59", x"EBD0", x"EB03", x"EB30", x"ED33", x"EF86", x"F167", x"F2DE", x"F2D6", x"F12B", x"F077", x"F1DA", x"F4D1", x"F953", x"FE5C", x"0143", x"01BC", x"00C2", x"FECB", x"FCF3", x"FCF7", x"FEAA", x"013C", x"0483", x"0769", x"08EF", x"09A1", x"09BA", x"08F4", x"0855", x"089C", x"0927", x"0A3E", x"0C0D", x"0D29", x"0CF5", x"0C55", x"0B1C", x"092D", x"07F9", x"0787", x"06CF", x"064F", x"064E", x"0579", x"040B", x"02DE", x"0115", x"FEA0", x"FD24", x"FC7C", x"FB96", x"FB04", x"FA40", x"F7C7", x"F4D6", x"F3CF", x"F4D5", x"F7F5", x"FD55", x"0279", x"04C4", x"049B", x"02C5", x"FF6E", x"FC76", x"FB77", x"FBC3", x"FCCD", x"FEC2", x"004A", x"0012", x"FEAA", x"FC5C", x"F931", x"F678", x"F534", x"F4BD", x"F4C2", x"F551", x"F5AF", x"F5A2", x"F5CD", x"F618", x"F5F9", x"F5B0", x"F52E", x"F437", x"F301", x"F1CE", x"F01A", x"EE6B", x"ED3D", x"ECBF", x"ED59", x"EFCF", x"F33F", x"F6A0", x"F988", x"FAF2", x"FA42", x"F941", x"FA0D", x"FCFD", x"0227", x"08E3", x"0E4F", x"104F", x"0F8E", x"0CD5", x"08B2", x"04FD", x"02FF", x"01E2", x"015F", x"01ED", x"0281", x"0212", x"017D", x"00CB", x"FFDE", x"FF93", x"0077", x"01BB", x"030E", x"04AD", x"05E6", x"06A9", x"0769", x"07F2", x"0824", x"088C", x"08F7", x"0926", x"0963", x"095B", x"0863", x"0757", x"064F", x"04DC", x"03F2", x"04B9", x"05FC", x"074E", x"08B7", x"0856", x"0550", x"026A", x"018E", x"0269", x"05D3", x"0B39", x"0EFE", x"0FF3", x"0FDD", x"0E8D", x"0BC5", x"09A9", x"0885", x"06DA", x"05A6", x"05B8", x"054F", x"03E8", x"02A8", x"00EB", x"FEB0", x"FD84", x"FD4E", x"FCFE", x"FCE6", x"FCDB", x"FBFB", x"FAF8", x"FA74", x"FA1A", x"FA9F", x"FC95", x"FEC2", x"00E2", x"0326", x"0449", x"0421", x"0414", x"03B5", x"026D", x"0223", x"0339", x"0412", x"0518", x"062F", x"04C2", x"013F", x"FEDC", x"FE30", x"FF25", x"0308", x"07F9", x"0A6B", x"0A8A", x"0979", x"0666", x"02AE", x"0097", x"FF9E", x"FF10", x"0005", x"0156", x"0132", x"0013", x"FE34", x"FB14", x"F81E", x"F676", x"F56B", x"F51F", x"F5BC", x"F5EA", x"F551", x"F4E4", x"F449", x"F3AA", x"F493", x"F6A1", x"F8D6", x"FBE2", x"FF8A", x"0212", x"03F1", x"0586", x"0518", x"0324", x"01C6", x"00D9", x"0000", x"006E", x"00D4", x"FF1B", x"FCD9", x"FC18", x"FCBD", x"FFDC", x"05F1", x"0C12", x"0FEF", x"1239", x"12C5", x"1181", x"10CA", x"1188", x"12B9", x"148C", x"170A", x"185D", x"17F1", x"167E", x"1397", x"0F8E", x"0C26", x"09B6", x"07DC", x"0749", x"07A3", x"07B7", x"07EA", x"088A", x"08D3", x"091A", x"0A08", x"0AAD", x"0AC3", x"0B0F", x"0ABE", x"0961", x"080F", x"06DA", x"04FE", x"03D8", x"0417", x"0467", x"04B6", x"050A", x"0328", x"FE7F", x"F999", x"F5E3", x"F424", x"F61A", x"FAF8", x"FEDD", x"003C", x"FF60", x"FBAF", x"F640", x"F210", x"EF78", x"EDF1", x"EE7B", x"F11E", x"F3FD", x"F6CB", x"F992", x"FB13", x"FB35", x"FB6F", x"FBD8", x"FC18", x"FCE1", x"FDFE", x"FEBC", x"FF8C", x"0098", x"0189", x"02D4", x"04D2", x"0718", x"09D9", x"0CF2", x"0F3E", x"10C9", x"1237", x"12DE", x"1298", x"12DA", x"136A", x"137F", x"145C", x"1571", x"145C", x"1146", x"0E59", x"0BAB", x"0A67", x"0C96", x"109E", x"132C", x"1460", x"148F", x"1295", x"0FD4", x"0E5C", x"0D41", x"0C34", x"0CDB", x"0EA9", x"0FFE", x"111F", x"11F1", x"116A", x"1074", x"103E", x"1022", x"0FF5", x"0FBE", x"0EC6", x"0CD4", x"0ABA", x"084D", x"0600", x"0506", x"050B", x"053E", x"0612", x"0670", x"0509", x"0358", x"0263", x"00F1", x"FFDB", x"00C6", x"0277", x"0461", x"07FA", x"0B25", x"0A9B", x"07AE", x"0455", x"00B4", x"FF42", x"0231", x"06BC", x"0A23", x"0D0C", x"0EAB", x"0E0B", x"0D30", x"0D88", x"0E15", x"0F84", x"12C2", x"1653", x"1924", x"1B85", x"1CCB", x"1CEA", x"1D28", x"1D90", x"1DD8", x"1E84", x"1F05", x"1E79", x"1D88", x"1C16", x"1971", x"1715", x"1606", x"1525", x"14B5", x"1591", x"15FE", x"158F", x"15EA", x"1634", x"1468", x"11F9", x"0FE8", x"0D1F", x"0B54", x"0C02", x"0C64", x"0AC7", x"08FA", x"076A", x"0645", x"0829", x"0D28", x"11B7", x"14BB", x"1647", x"1521", x"120F", x"0F83", x"0DB7", x"0C45", x"0C25", x"0C91", x"0C0D", x"0AFF", x"0974", x"06BE", x"03E5", x"01E1", x"000C", x"FF12", x"FFB3", x"00C0", x"0160", x"0238", x"0248", x"0112", x"004D", x"0047", x"FFD0", x"FF9F", x"FFC3", x"FE9E", x"FCB4", x"FB91", x"FA44", x"F8B6", x"F8AE", x"FA00", x"FBC0", x"FF2C", x"03A9", x"0635", x"06AB", x"064C", x"051B", x"04CA", x"07DC", x"0D1F", x"11F9", x"15C4", x"174E", x"154A", x"1183", x"0DE5", x"0A68", x"07D9", x"0756", x"07B0", x"0843", x"09AC", x"0AEF", x"0B1B", x"0B09", x"0AF2", x"0A3B", x"0A3B", x"0B60", x"0C95", x"0DCB", x"0F73", x"1070", x"10EA", x"1215", x"1346", x"13DD", x"14A8", x"14EE", x"139D", x"122D", x"1149", x"0FBA", x"0E54", x"0E1F", x"0DB2", x"0D3A", x"0EAC", x"106F", x"1046", x"0F27", x"0D66", x"0A70", x"090B", x"0B7D", x"0F5D", x"12D8", x"1619", x"1734", x"1504", x"1210", x"0F29", x"0B8E", x"087A", x"0753", x"0676", x"05C1", x"05C3", x"053E", x"0385", x"024A", x"01A5", x"0123", x"0182", x"0256", x"023F", x"01AE", x"012A", x"003A", x"FFC0", x"0089", x"0199", x"02BD", x"0467", x"052D", x"0499", x"043B", x"03B7", x"0224", x"0135", x"0134", x"00E1", x"01C1", x"04E0", x"0771", x"07B2", x"06B8", x"03F5", x"0005", x"FEEE", x"01C8", x"05E6", x"0A67", x"0EAA", x"100E", x"0EC4", x"0D13", x"0AF5", x"083C", x"06B2", x"05FB", x"04CD", x"03D3", x"02F7", x"011E", x"FF16", x"FDB8", x"FC11", x"FA8B", x"FA21", x"F983", x"F864", x"F7EE", x"F754", x"F651", x"F6C9", x"F8DF", x"FAFB", x"FE09", x"01CD", x"042D", x"05C3", x"07FD", x"08F8", x"07C7", x"063E", x"03A7", x"FFA9", x"FD7D", x"FDDA", x"FDA9", x"FC94", x"FB6B", x"F8CB", x"F667", x"F806", x"FCF6", x"027D", x"0879", x"0D9F", x"0FB3", x"102F", x"10F1", x"10E6", x"1038", x"1042", x"0FEE", x"0E78", x"0D42", x"0BC6", x"08FD", x"060B", x"0396", x"00EF", x"FF57", x"FFA7", x"0090", x"017C", x"02FA", x"0402", x"0473", x"0591", x"0731", x"0861", x"09D5", x"0B24", x"0B4C", x"0B06", x"0ACE", x"0999", x"07FE", x"06EA", x"0578", x"040A", x"0416", x"0486", x"0380", x"01A3", x"FE92", x"F9E1", x"F66C", x"F680", x"F8CE", x"FC23", x"FFFB", x"018D", x"FF8D", x"FC3C", x"F8A5", x"F495", x"F20B", x"F1C9", x"F205", x"F2F3", x"F548", x"F73B", x"F806", x"F8F8", x"F96F", x"F8E3", x"F922", x"FA57", x"FAF2", x"FB64", x"FC51", x"FC9E", x"FD06", x"FEFF", x"016E", x"03C1", x"06AB", x"092A", x"0A4A", x"0B82", x"0C89", x"0BFF", x"0AE3", x"099B", x"06A5", x"03C9", x"034A", x"035B", x"028E", x"01E9", x"FFBC", x"FB40", x"F897", x"F9A8", x"FBE1", x"FEE9", x"02CE", x"042F", x"028A", x"0140", x"0000", x"FD4B", x"FB8C", x"FB6E", x"FABD", x"FA52", x"FB3E", x"FAEB", x"F8BF", x"F725", x"F5BC", x"F3F1", x"F32C", x"F2E5", x"F10C", x"EE7D", x"EC7E", x"EA95", x"E967", x"E994", x"E9CF", x"E9B4", x"E9D1", x"E982", x"E8E1", x"E8DE", x"E8D6", x"E87D", x"E957", x"EAA5", x"EBC7", x"EE91", x"F2F0", x"F60C", x"F786", x"F773", x"F3C9", x"EE4E", x"EBCA", x"EC68", x"EE8F", x"F2E8", x"F791", x"F93D", x"F99E", x"FAF8", x"FBDE", x"FCB2", x"FF6A", x"0259", x"0445", x"06EB", x"098A", x"0A24", x"09F7", x"098F", x"0784", x"0517", x"03C4", x"01FB", x"FFC9", x"FE6D", x"FCDA", x"FAC1", x"FA22", x"FA5F", x"FA39", x"FAEF", x"FC06", x"FBD5", x"FBD1", x"FCF2", x"FCEE", x"FBF5", x"FB1B", x"F864", x"F422", x"F237", x"F262", x"F22A", x"F295", x"F2AD", x"EFB2", x"EC64", x"ECBD", x"EEF4", x"F18C", x"F59F", x"F880", x"F7FA", x"F724", x"F757", x"F640", x"F4BD", x"F45B", x"F321", x"F106", x"F034", x"EF7C", x"ED39", x"EAFB", x"E93D", x"E6FC", x"E5A8", x"E5FD", x"E64A", x"E62C", x"E66D", x"E64C", x"E5D6", x"E602", x"E676", x"E6B0", x"E73E", x"E7BB", x"E7B4", x"E7F0", x"E82A", x"E812", x"E8C1", x"EA30", x"EB3D", x"ECF1", x"F03C", x"F343", x"F590", x"F768", x"F690", x"F286", x"EF18", x"EE1A", x"EED9", x"F240", x"F795", x"FAB6", x"FB0A", x"FAA8", x"F922", x"F655", x"F4CB", x"F47B", x"F393", x"F36F", x"F4AC", x"F525", x"F4F8", x"F55C", x"F53D", x"F46D", x"F4B5", x"F596", x"F5B6", x"F62F", x"F6FF", x"F725", x"F78D", x"F8A3", x"F91F", x"F918", x"F946", x"F892", x"F754", x"F6DF", x"F655", x"F539", x"F4E1", x"F441", x"F230", x"F11D", x"F211", x"F33C", x"F4CA", x"F726", x"F705", x"F4A5", x"F44A", x"F64C", x"F8EA", x"FD39", x"01ED", x"0328", x"01CF", x"00F7", x"FEF6", x"FB57", x"F8D4", x"F6DE", x"F3EF", x"F20B", x"F1D2", x"F0B0", x"EEFC", x"EEB3", x"EEF0", x"EF6D", x"F12C", x"F2F8", x"F30F", x"F242", x"F164", x"F035", x"EF52", x"EF05", x"EEC2", x"EEE3", x"EF88", x"F077", x"F1C6", x"F321", x"F36A", x"F36D", x"F3BB", x"F333", x"F267", x"F331", x"F4A3", x"F587", x"F6B9", x"F6CB", x"F367", x"EF22", x"ED76", x"ED9C", x"EFC1", x"F492", x"F8E8", x"FA28", x"FA97", x"FB18", x"FA0A", x"F8A4", x"F825", x"F6C5", x"F4B6", x"F3F4", x"F38B", x"F268", x"F189", x"F0D9", x"EF3B", x"EDC3", x"ECCC", x"EB5A", x"E9FB", x"E957", x"E8C4", x"E8BC", x"E9E6", x"EB3E", x"EC9A", x"EEBC", x"F060", x"F122", x"F255", x"F3A9", x"F403", x"F4CE", x"F5B2", x"F475", x"F27E", x"F22B", x"F257", x"F2F3", x"F534", x"F6BB", x"F55D", x"F479", x"F5F9", x"F870", x"FC58", x"0204", x"05DB", x"06BE", x"0786", x"0818", x"0720", x"0644", x"0620", x"04DD", x"0363", x"02FA", x"0236", x"0050", x"FE88", x"FCBD", x"FA99", x"F95F", x"F92D", x"F947", x"F9D1", x"FB08", x"FC44", x"FDAF", x"FF22", x"0034", x"010B", x"01F7", x"0244", x"0246", x"021D", x"0114", x"FF68", x"FE50", x"FCE8", x"FAA3", x"F8FE", x"F829", x"F708", x"F681", x"F65D", x"F3EC", x"EF69", x"EBAE", x"E964", x"E8BB", x"EB45", x"EF8F", x"F245", x"F38D", x"F46A", x"F3DA", x"F265", x"F1D5", x"F188", x"F0C5", x"F0BE", x"F157", x"F16C", x"F17C", x"F1FE", x"F219", x"F203", x"F22F", x"F200", x"F1A0", x"F1F1", x"F2EC", x"F4B5", x"F7B7", x"FB21", x"FE64", x"01FF", x"055D", x"07B2", x"09B0", x"0AF2", x"0A86", x"099C", x"092F", x"07E3", x"0625", x"05CA", x"0618", x"0661", x"0809", x"09A7", x"0872", x"05E9", x"0493", x"0418", x"0501", x"08CF", x"0CDD", x"0EC0", x"1005", x"115F", x"1160", x"10D5", x"10FA", x"104E", x"0EB2", x"0DBC", x"0CF6", x"0B2E", x"094F", x"07E2", x"064D", x"052E", x"04C3", x"0447", x"0346", x"0244", x"013C", x"0067", x"FFBF", x"FEDF", x"FDC4", x"FCCF", x"FBD0", x"FB10", x"FB05", x"FAC9", x"FA12", x"F9FD", x"FA4E", x"FA24", x"FA6B", x"FBC7", x"FCD6", x"FDC2", x"FF02", x"FEA2", x"FB76", x"F7F0", x"F593", x"F462", x"F5AB", x"F993", x"FD8A", x"00A2", x"041B", x"079D", x"0A5D", x"0D0C", x"0F98", x"10EC", x"115F", x"1180", x"10EF", x"0F9A", x"0E32", x"0CD1", x"0BA9", x"0ACE", x"0A03", x"0930", x"08BA", x"0838", x"07F4", x"085A", x"08CA", x"08FA", x"09F3", x"0B7B", x"0CA2", x"0DE9", x"0F75", x"0FF2", x"0FE2", x"108A", x"1075", x"0E96", x"0C78", x"0A61", x"07B2", x"061E", x"061A", x"0508", x"025F", x"006B", x"FF58", x"FF0A", x"011F", x"04B8", x"06F5", x"07F4", x"08E0", x"08CF", x"079D", x"06A1", x"053B", x"02C3", x"0074", x"FEDF", x"FD31", x"FBC2", x"FAFA", x"FA17", x"F91F", x"F890", x"F813", x"F764", x"F70E", x"F6C3", x"F64E", x"F600", x"F5BF", x"F52F", x"F4F5", x"F536", x"F592", x"F680", x"F7F9", x"F94F", x"FAD8", x"FD0C", x"FF00", x"005B", x"01D6", x"02EA", x"031A", x"0345", x"02E7", x"007A", x"FCD8", x"F9BA", x"F794", x"F761", x"FA29", x"FE60", x"01FD", x"04EF", x"06FA", x"0762", x"070D", x"06C6", x"0629", x"053C", x"04AA", x"03E5", x"02F6", x"0286", x"0286", x"02B2", x"036E", x"0432", x"049A", x"052A", x"0614", x"06EE", x"083C", x"09FB", x"0B2D", x"0C1C", x"0D54", x"0E06", x"0E2A", x"0E84", x"0E25", x"0C9F", x"0B7E", x"0AC6", x"0941", x"07F6", x"07B5", x"073D", x"0752", x"0937", x"0AE9", x"0A9D", x"09FB", x"097D", x"08BB", x"099E", x"0CC7", x"0F75", x"10C1", x"11FC", x"1254", x"1142", x"1076", x"0FAB", x"0D9F", x"0B53", x"09E0", x"084B", x"06ED", x"0688", x"065F", x"05FF", x"0651", x"06C8", x"0690", x"05CF", x"0479", x"021F", x"FF97", x"FD6F", x"FB91", x"FA7A", x"FA84", x"FB0E", x"FC43", x"FDEA", x"FF09", x"FF87", x"0056", x"00E1", x"00E5", x"0161", x"021A", x"022E", x"02B1", x"03AE", x"031D", x"00DF", x"FE56", x"FBCA", x"F9E8", x"FA97", x"FD30", x"FF9F", x"01D1", x"03E9", x"051E", x"05CD", x"06B1", x"070A", x"064B", x"052A", x"036C", x"0116", x"FEE2", x"FD0B", x"FB59", x"FA3F", x"F9B6", x"F944", x"F953", x"FA0E", x"FAE1", x"FC05", x"FDC3", x"FF40", x"009B", x"028A", x"0470", x"0595", x"06C2", x"0762", x"06BC", x"0628", x"0690", x"068E", x"060B", x"0600", x"057B", x"0495", x"0564", x"0784", x"08A2", x"0923", x"09BA", x"09D3", x"0A51", x"0CF9", x"1052", x"12A0", x"148A", x"1634", x"16AF", x"170C", x"17F2", x"1825", x"1772", x"1676", x"14B3", x"11DA", x"0EFE", x"0C47", x"097A", x"0761", x"062C", x"055B", x"0512", x"05AC", x"0661", x"0740", x"0892", x"09BF", x"0ABD", x"0C22", x"0D9B", x"0EDC", x"1061", x"118B", x"11D5", x"1201", x"1260", x"11F4", x"1126", x"106E", x"0EF3", x"0CF5", x"0BE0", x"0A93", x"07D8", x"049C", x"0198", x"FEA4", x"FD8E", x"FF56", x"023E", x"0508", x"07FC", x"09FB", x"0A5A", x"0A57", x"0A1D", x"08D4", x"0739", x"05D0", x"03BC", x"01AE", x"008F", x"FFF3", x"FFCF", x"0100", x"02C1", x"0460", x"067C", x"08B5", x"0A61", x"0C41", x"0EB5", x"10EC", x"1310", x"1569", x"16A8", x"16EB", x"16E0", x"15EB", x"1416", x"12EA", x"11EA", x"1072", x"0F8F", x"0F6A", x"0EC1", x"0ED8", x"103A", x"10D4", x"0FF5", x"0F31", x"0E1B", x"0D0A", x"0E3B", x"117A", x"1446", x"16C2", x"1901", x"1985", x"18C9", x"1836", x"16BD", x"13DF", x"10FC", x"0DC5", x"09A4", x"05F2", x"0312", x"FFE3", x"FD65", x"FC30", x"FB55", x"FAC6", x"FB2C", x"FB1F", x"FA2B", x"F952", x"F84F", x"F6F1", x"F66F", x"F6B5", x"F6E8", x"F7DD", x"F978", x"FA75", x"FB8C", x"FD7A", x"FECE", x"FF68", x"0075", x"00A8", x"FFC0", x"FFC8", x"004C", x"FF1C", x"FCF5", x"FAC1", x"F7DB", x"F622", x"F80D", x"FC0D", x"0041", x"0527", x"09D7", x"0D2E", x"10AB", x"14C6", x"17B6", x"1953", x"1A24", x"194F", x"1721", x"1538", x"1380", x"11B7", x"10BF", x"109C", x"1056", x"1054", x"1047", x"0F60", x"0DF6", x"0CBC", x"0B8D", x"0AF8", x"0B7B", x"0C47", x"0D50", x"0ED6", x"0FCB", x"0FE3", x"103E", x"1096", x"1026", x"0FD4", x"0F5A", x"0D6B", x"0B16", x"0A03", x"0908", x"0787", x"065F", x"0507", x"0320", x"02DB", x"050B", x"0805", x"0B1B", x"0E25", x"0FB8", x"0F93", x"0F13", x"0E2B", x"0C8B", x"0AD8", x"08FB", x"0658", x"0349", x"006B", x"FD81", x"FB21", x"F9AC", x"F889", x"F76D", x"F688", x"F57A", x"F44B", x"F3C2", x"F3AD", x"F3BE", x"F473", x"F5B7", x"F6F4", x"F8EA", x"FB8A", x"FDB8", x"FF90", x"01F0", x"040D", x"0562", x"06BB", x"074F", x"0614", x"0460", x"035D", x"018D", x"FEC0", x"FC14", x"F973", x"F725", x"F759", x"FA76", x"FE3F", x"020B", x"05F5", x"08EB", x"0A95", x"0C2A", x"0D7B", x"0DA9", x"0D2E", x"0C6B", x"0A84", x"079D", x"0492", x"019E", x"FF31", x"FE23", x"FE52", x"FED1", x"FF3F", x"FF65", x"FF1A", x"FEF4", x"FF5F", x"004E", x"0160", x"0236", x"0277", x"0258", x"0201", x"012A", x"003F", x"FF72", x"FE5F", x"FD2C", x"FCC2", x"FCC8", x"FD39", x"FEFC", x"01C6", x"03BC", x"0492", x"04C8", x"0412", x"0357", x"0450", x"0683", x"0866", x"09F7", x"0B31", x"0B32", x"0A8A", x"0A08", x"090D", x"0799", x"0639", x"04A4", x"02A1", x"00E5", x"FF8D", x"FE57", x"FDEB", x"FE08", x"FDE5", x"FDB8", x"FD80", x"FC84", x"FAF6", x"F9AB", x"F82C", x"F6C7", x"F645", x"F62D", x"F5E3", x"F613", x"F669", x"F622", x"F631", x"F6ED", x"F71F", x"F709", x"F746", x"F6C8", x"F5B2", x"F5BF", x"F60A", x"F4D6", x"F2D2", x"F074", x"ED4A", x"EB65", x"ECA0", x"EF63", x"F229", x"F533", x"F789", x"F87B", x"F970", x"FAFC", x"FBF1", x"FC50", x"FC6F", x"FB42", x"F8DC", x"F643", x"F393", x"F0DC", x"EF2D", x"EE7B", x"EE3E", x"EE90", x"EF2F", x"EF54", x"EF20", x"EEF4", x"EEB2", x"EE9B", x"EEC0", x"EEEB", x"EF31", x"EFC9", x"F03F", x"F0C2", x"F1D4", x"F2FD", x"F451", x"F665", x"F876", x"F995", x"FACC", x"FC92", x"FDDC", x"FEA5", x"FF49", x"FEC3", x"FD58", x"FD43", x"FEE7", x"013B", x"041C", x"0708", x"0891", x"08F3", x"0934", x"093A", x"08D1", x"0876", x"07A2", x"05B9", x"0317", x"003C", x"FD70", x"FB7F", x"FAC7", x"FA9A", x"FA9E", x"FA8A", x"F9F5", x"F938", x"F8F4", x"F920", x"F99A", x"FA82", x"FB1D", x"FB6B", x"FC08", x"FCB4", x"FCE4", x"FCDF", x"FCDB", x"FC01", x"FAF6", x"FA56", x"F915", x"F6CA", x"F4CC", x"F310", x"F075", x"ED4A", x"EA3A", x"E6BB", x"E3F5", x"E42D", x"E71B", x"EACE", x"EEB9", x"F25B", x"F44A", x"F4CC", x"F4F0", x"F482", x"F2DD", x"F0CF", x"EE85", x"EB60", x"E7B9", x"E481", x"E235", x"E142", x"E236", x"E4A7", x"E75A", x"E9CA", x"EBBA", x"ED5C", x"EF0A", x"F109", x"F356", x"F568", x"F6DF", x"F7CC", x"F886", x"F8F0", x"F8ED", x"F8F9", x"F8E3", x"F83C", x"F789", x"F719", x"F657", x"F564", x"F599", x"F650", x"F635", x"F58E", x"F47D", x"F2BC", x"F1C1", x"F377", x"F6CF", x"FA47", x"FDDE", x"0105", x"02C7", x"03B8", x"0475", x"0420", x"029F", x"00B1", x"FE1B", x"FACF", x"F782", x"F494", x"F24C", x"F13A", x"F10D", x"F11B", x"F169", x"F1BA", x"F187", x"F163", x"F161", x"F0CC", x"F003", x"EF9C", x"EF04", x"EE53", x"EE4E", x"EE39", x"EDA1", x"ED85", x"EDBD", x"ED59", x"ED0B", x"ECF4", x"EBE2", x"EAAF", x"EAE7", x"EB52", x"EB1D", x"EAED", x"EA26", x"E874", x"E841", x"EABE", x"EE6D", x"F2BA", x"F78D", x"FB16", x"FD37", x"FF47", x"0130", x"0278", x"03D3", x"0494", x"03BB", x"0210", x"0028", x"FDDF", x"FC76", x"FC53", x"FC27", x"FBFA", x"FC83", x"FCFD", x"FD0D", x"FDDA", x"FE94", x"FE85", x"FEE0", x"FFD5", x"0079", x"0168", x"02E9", x"03AC", x"03E4", x"046E", x"043D", x"034B", x"02A3", x"015F", x"FED6", x"FCDD", x"FBA1", x"F9E9", x"F85B", x"F718", x"F48D", x"F1D2", x"F174", x"F2FD", x"F5C1", x"F9F5", x"FDEB", x"FFAA", x"003A", x"0051", x"FF59", x"FE45", x"FD99", x"FBEE", x"F920", x"F61E", x"F2B7", x"EF37", x"ED1B", x"EBBB", x"E9F0", x"E83B", x"E696", x"E466", x"E2E8", x"E2D1", x"E34D", x"E473", x"E66D", x"E81B", x"E991", x"EBCA", x"EE08", x"EFEF", x"F23B", x"F42A", x"F4F5", x"F631", x"F7CE", x"F81C", x"F7AB", x"F78B", x"F658", x"F441", x"F2C5", x"F0A7", x"ED10", x"EA90", x"EA8D", x"EC03", x"EF64", x"F443", x"F806", x"FA0A", x"FBD4", x"FD45", x"FE27", x"FF7D", x"008F", x"FFFD", x"FE5D", x"FC39", x"F95C", x"F712", x"F641", x"F5F0", x"F5F1", x"F6A0", x"F737", x"F79F", x"F8DA", x"FA9A", x"FC0F", x"FDEE", x"FFD3", x"00E3", x"01DC", x"0333", x"03A7", x"0379", x"0355", x"0262", x"00AA", x"FFE8", x"FF90", x"FE7B", x"FE06", x"FEC9", x"FF74", x"000E", x"010C", x"00A8", x"FE91", x"FD4B", x"FDCC", x"FF4C", x"021B", x"05B4", x"086F", x"0A12", x"0B84", x"0C50", x"0C0B", x"0B16", x"0953", x"06A4", x"03A6", x"009A", x"FDC2", x"FBCB", x"FAA2", x"F97E", x"F86A", x"F71E", x"F530", x"F38E", x"F305", x"F2F3", x"F320", x"F3E3", x"F465", x"F465", x"F52D", x"F68E", x"F79F", x"F8E5", x"FA8F", x"FB4B", x"FBE0", x"FD3C", x"FDE3", x"FD42", x"FCD9", x"FC90", x"FB72", x"FA9F", x"F9C5", x"F6FF", x"F33D", x"F114", x"F077", x"F1A3", x"F516", x"F912", x"FB80", x"FD1D", x"FE3D", x"FE56", x"FE97", x"FF6D", x"FF43", x"FE23", x"FCD6", x"FAAB", x"F843", x"F768", x"F748", x"F699", x"F682", x"F702", x"F70D", x"F7B2", x"F99B", x"FA92", x"FA7C", x"FA9A", x"FA57", x"F978", x"F9D8", x"FB06", x"FBE2", x"FD84", x"FFF9", x"01DE", x"03B1", x"0611", x"0750", x"07AC", x"08DF", x"0A33", x"0B05", x"0C58", x"0CE6", x"0B52", x"095C", x"08E7", x"097C", x"0BDF", x"1027", x"13E3", x"1605", x"1769", x"17A0", x"168E", x"1591", x"146B", x"11DE", x"0EE6", x"0BD4", x"080F", x"04E4", x"033C", x"01B0", x"FFF4", x"FED0", x"FD8C", x"FC0B", x"FBE1", x"FCBA", x"FDA8", x"FF4E", x"016B", x"02E6", x"049D", x"06F4", x"08E3", x"0AAD", x"0CA8", x"0D45", x"0CC3", x"0CF3", x"0CF0", x"0BCB", x"0AF4", x"09DA", x"0710", x"0449", x"0278", x"FF4D", x"FB06", x"F838", x"F694", x"F64A", x"F94D", x"FE00", x"011E", x"030A", x"0459", x"040D", x"036C", x"03F7", x"0405", x"02AA", x"0177", x"000D", x"FE2E", x"FDA9", x"FE7A", x"FEF0", x"FF7A", x"00AC", x"01A0", x"02A0", x"04B5", x"06B1", x"07E5", x"0925", x"09DF", x"09C5", x"09ED", x"0A60", x"0A61", x"0A8C", x"0B13", x"0AAB", x"0A59", x"0B0F", x"0B95", x"0B70", x"0C04", x"0CA5", x"0CCA", x"0DB8", x"0F27", x"0EB3", x"0CEB", x"0BB5", x"0B47", x"0C11", x"0F27", x"1309", x"15A5", x"171F", x"17E4", x"172F", x"1587", x"134E", x"1043", x"0C62", x"0878", x"0486", x"00BD", x"FDBA", x"FB50", x"F967", x"F80C", x"F6EB", x"F5C1", x"F54B", x"F5B6", x"F6A5", x"F839", x"FA10", x"FAE6", x"FB28", x"FB94", x"FBD8", x"FC0A", x"FCF5", x"FD82", x"FCE9", x"FC8F", x"FCB1", x"FBF0", x"FB0C", x"FAF0", x"FABD", x"FAA3", x"FC17", x"FD8E", x"FCE2", x"FB64", x"FA68", x"F9E9", x"FB63", x"FFB5", x"046B", x"07F0", x"0ADA", x"0CB5", x"0D56", x"0E4F", x"0FF6", x"10FC", x"11F2", x"12F6", x"12DC", x"123F", x"121C", x"1166", x"0FA5", x"0E57", x"0D18", x"0B83", x"0B17", x"0BB7", x"0B65", x"0A92", x"0A16", x"08FE", x"07E1", x"0852", x"096B", x"0A3A", x"0BE8", x"0DD6", x"0EAF", x"0F7C", x"106E", x"0FEC", x"0EEA", x"0ED8", x"0EE0", x"0EBE", x"0F7F", x"0F5C", x"0D0B", x"0AB1", x"09B2", x"09DE", x"0C2E", x"10A2", x"145D", x"1672", x"178F", x"170B", x"14E7", x"12AF", x"1020", x"0CA2", x"0952", x"0641", x"02B0", x"FFAF", x"FD98", x"FB2C", x"F8A7", x"F71B", x"F5B5", x"F4AE", x"F546", x"F690", x"F76B", x"F8A8", x"FA03", x"FAA3", x"FB81", x"FD09", x"FE2F", x"FF76", x"0129", x"01F3", x"0232", x"0325", x"03AF", x"035A", x"037A", x"0341", x"01B6", x"00F8", x"0115", x"FF8E", x"FD44", x"FBE2", x"FAC6", x"FB3B", x"FFA6", x"05B3", x"0A69", x"0E3C", x"10AC", x"106F", x"1016", x"1110", x"111B", x"1010", x"0F25", x"0CCC", x"08FA", x"0657", x"0450", x"0146", x"FF10", x"FE38", x"FD4A", x"FD53", x"FF51", x"00C3", x"0137", x"0223", x"02DD", x"02E5", x"0401", x"0586", x"05F8", x"065E", x"06CF", x"05FD", x"0549", x"0594", x"0538", x"042F", x"0411", x"03C8", x"035B", x"04F7", x"075D", x"07E3", x"0770", x"073E", x"06AA", x"07C1", x"0C26", x"1163", x"1568", x"18B1", x"1A4D", x"198B", x"1832", x"16CD", x"1463", x"11BC", x"0F7F", x"0CAC", x"09E7", x"07F6", x"061C", x"0436", x"031C", x"01FF", x"00BC", x"0094", x"0148", x"0216", x"03A3", x"053E", x"0575", x"0537", x"0549", x"04CF", x"04B9", x"05C0", x"05FD", x"052C", x"052B", x"0522", x"0406", x"036D", x"032C", x"016E", x"0015", x"00B1", x"0094", x"FEE4", x"FD62", x"FB76", x"F973", x"FAB4", x"FF34", x"03DB", x"081F", x"0BB1", x"0C9B", x"0BE5", x"0C05", x"0C35", x"0BEF", x"0C73", x"0C64", x"0A87", x"08AB", x"0727", x"0492", x"0221", x"00DA", x"FF39", x"FE0E", x"FF0E", x"0082", x"00E0", x"014A", x"0107", x"FF28", x"FDE7", x"FE56", x"FEE7", x"004B", x"031B", x"0579", x"0726", x"0993", x"0B82", x"0BE9", x"0C70", x"0D33", x"0D23", x"0DCF", x"0F7F", x"0FAE", x"0E15", x"0C6B", x"0AB9", x"09FA", x"0C68", x"1117", x"15C9", x"19F3", x"1CF1", x"1D92", x"1CD6", x"1BEE", x"1A8F", x"1958", x"18C4", x"177D", x"1555", x"1323", x"1056", x"0CE3", x"0A30", x"07DA", x"0520", x"0361", x"02D8", x"0245", x"023B", x"0350", x"0419", x"04DC", x"06E0", x"08FC", x"0AB0", x"0CFA", x"0ED2", x"0EF4", x"0F0D", x"0F8C", x"0ED6", x"0DEA", x"0D5C", x"0B17", x"0795", x"0570", x"035C", x"FFE9", x"FCC6", x"F9B2", x"F5DF", x"F457", x"F6E3", x"FAED", x"FF1D", x"035E", x"050D", x"03F4", x"033A", x"0349", x"030F", x"03D5", x"04DB", x"03A6", x"0174", x"FFE7", x"FDA7", x"FB29", x"FA3E", x"F9A4", x"F8C1", x"F9AE", x"FBE3", x"FD2A", x"FE68", x"FFDA", x"0005", x"0001", x"015A", x"0293", x"035A", x"04DA", x"05D9", x"05D7", x"0693", x"07CF", x"080D", x"0863", x"08EE", x"082D", x"077A", x"084C", x"08DA", x"082A", x"0764", x"0620", x"0485", x"0565", x"0929", x"0DD0", x"12AB", x"16EC", x"18D6", x"18CA", x"1818", x"16A4", x"14DC", x"138B", x"11A8", x"0EBA", x"0BDC", x"08CF", x"059D", x"03B1", x"029B", x"00CE", x"FF3D", x"FE77", x"FD85", x"FD43", x"FE94", x"FF64", x"FF0A", x"FEEF", x"FE67", x"FD26", x"FD47", x"FE59", x"FE21", x"FDD1", x"FE42", x"FDD6", x"FD2F", x"FE0A", x"FE4F", x"FD3B", x"FD81", x"FEE8", x"FF42", x"FF62", x"FF55", x"FD2A", x"FABA", x"FB04", x"FD39", x"0028", x"03EE", x"0688", x"0638", x"04D3", x"03A1", x"0274", x"02C0", x"04CF", x"066F", x"075F", x"084C", x"085F", x"07AD", x"07EF", x"086A", x"082E", x"0889", x"099C", x"09CA", x"0987", x"092E", x"0793", x"0521", x"03AB", x"02C4", x"0234", x"02DD", x"0426", x"04F0", x"05E3", x"0720", x"0780", x"075A", x"0759", x"06A7", x"059F", x"0570", x"0589", x"04B5", x"0348", x"014F", x"FF00", x"FDC3", x"FEC0", x"0167", x"04BC", x"07CA", x"095E", x"08FA", x"06D1", x"0354", x"FFCC", x"FD1C", x"FAF6", x"F8D9", x"F6B8", x"F3B1", x"EFE1", x"ECCB", x"EAFC", x"E98B", x"E8D7", x"E8F2", x"E8EB", x"E8C6", x"E9A2", x"EAB5", x"EB73", x"EC8E", x"EE10", x"EF14", x"F08E", x"F2D6", x"F4B5", x"F601", x"F7AE", x"F8DA", x"F92A", x"F9B7", x"FA26", x"F920", x"F7E4", x"F76E", x"F68B", x"F4D3", x"F31B", x"F0C9", x"EDED", x"ED1A", x"EF3F", x"F2B9", x"F6BB", x"FA86", x"FC61", x"FC3C", x"FBEB", x"FBD2", x"FBE9", x"FCB9", x"FD8F", x"FD0B", x"FB81", x"F997", x"F730", x"F53A", x"F4BC", x"F4D3", x"F549", x"F6B8", x"F883", x"F991", x"FA9E", x"FBBA", x"FC32", x"FCB5", x"FDC8", x"FE6D", x"FE4F", x"FE30", x"FD77", x"FC16", x"FAED", x"F9D7", x"F80A", x"F658", x"F503", x"F3A4", x"F322", x"F47D", x"F627", x"F754", x"F86F", x"F951", x"F9FD", x"FC6F", x"00FC", x"05F4", x"0A8A", x"0E68", x"1054", x"100D", x"0E81", x"0BFC", x"08D0", x"05C6", x"02CF", x"FF97", x"FC1C", x"F843", x"F478", x"F1AA", x"EFBA", x"EE17", x"ED35", x"ED18", x"ED29", x"EDF2", x"EFF8", x"F1D9", x"F34D", x"F4FF", x"F62A", x"F666", x"F6E5", x"F770", x"F6F7", x"F678", x"F683", x"F5C1", x"F492", x"F3ED", x"F27C", x"F020", x"EF26", x"EF51", x"EEDF", x"EE4C", x"ED71", x"EADE", x"E81E", x"E801", x"E9C3", x"EC4D", x"EFD2", x"F2FE", x"F417", x"F43D", x"F450", x"F3B8", x"F33D", x"F383", x"F363", x"F264", x"F113", x"EEF9", x"EC36", x"EA46", x"E927", x"E858", x"E8C3", x"EA40", x"EB74", x"EC42", x"ED25", x"ED15", x"EC93", x"ECE6", x"EDBF", x"EEAD", x"F077", x"F2F5", x"F555", x"F811", x"FB18", x"FD25", x"FE67", x"FF6F", x"FFB5", x"FFBC", x"00D9", x"0241", x"029B", x"0223", x"00DE", x"FE9F", x"FD54", x"FEAA", x"01A1", x"0502", x"0879", x"0ABF", x"0AFD", x"09E9", x"083D", x"05E6", x"0397", x"01C7", x"FFF4", x"FDC4", x"FB4E", x"F860", x"F599", x"F37B", x"F1C7", x"F054", x"EF95", x"EF1C", x"EEDB", x"EF70", x"F0F4", x"F2C3", x"F547", x"F891", x"FBAB", x"FE9F", x"01DA", x"04B7", x"06F4", x"0954", x"0B1B", x"0B5F", x"0AE1", x"096B", x"0623", x"0272", x"FFC7", x"FCD6", x"F924", x"F59C", x"F17D", x"ECC8", x"EA7E", x"EBAC", x"EE1C", x"F146", x"F508", x"F75C", x"F81B", x"F940", x"FA8D", x"FB06", x"FBB3", x"FC98", x"FC38", x"FB0A", x"F9B2", x"F779", x"F4FD", x"F3AC", x"F306", x"F2D6", x"F403", x"F58F", x"F64D", x"F6E9", x"F770", x"F71A", x"F719", x"F803", x"F8A1", x"F916", x"FA14", x"FAB6", x"FB18", x"FC6C", x"FDED", x"FEAD", x"FFB3", x"005B", x"FFB6", x"FFB0", x"0110", x"01EE", x"0240", x"02A7", x"01BF", x"0010", x"00E8", x"03DC", x"06D5", x"0A38", x"0D7E", x"0E6E", x"0DFA", x"0D69", x"0B7A", x"07FF", x"04B0", x"013C", x"FD47", x"FA42", x"F7E2", x"F528", x"F301", x"F154", x"EF04", x"ED0D", x"EC2F", x"EB54", x"EACB", x"EB62", x"EBB5", x"EB71", x"EC01", x"EC9B", x"EC6B", x"ECBB", x"ED7A", x"ED78", x"EE1D", x"EFD1", x"F0C0", x"F122", x"F1B7", x"F0D4", x"EEF2", x"EEE1", x"EFFA", x"F094", x"F189", x"F1EF", x"EFE2", x"EDEA", x"EED2", x"F0FE", x"F3B1", x"F771", x"FA0C", x"FA28", x"FA13", x"FA4E", x"F9CE", x"F9CD", x"FAF9", x"FBCF", x"FC6D", x"FD9B", x"FE0B", x"FD9C", x"FD8B", x"FD24", x"FC21", x"FBDB", x"FC1F", x"FBC0", x"FB79", x"FB15", x"F97A", x"F799", x"F686", x"F59E", x"F533", x"F63C", x"F7A5", x"F924", x"FBA5", x"FE5B", x"004F", x"028D", x"0471", x"049F", x"0495", x"05BA", x"0693", x"0724", x"0807", x"072C", x"0433", x"0260", x"02CC", x"0410", x"0690", x"09C1", x"0AEE", x"0A09", x"0904", x"0752", x"0474", x"01FD", x"FFF0", x"FD6A", x"FB6C", x"FA41", x"F8C6", x"F706", x"F59E", x"F3B9", x"F179", x"EFF1", x"EEEF", x"EE2C", x"EE55", x"EF43", x"F028", x"F187", x"F345", x"F4B1", x"F610", x"F7A5", x"F8C0", x"F997", x"FAA2", x"FB49", x"FB93", x"FC83", x"FD01", x"FC5F", x"FC08", x"FC59", x"FC1B", x"FBD6", x"FBCC", x"FA2F", x"F790", x"F731", x"F925", x"FBE1", x"FFBB", x"03EA", x"0600", x"06AB", x"07B7", x"07FE", x"06C2", x"0588", x"0450", x"0238", x"003C", x"FEBD", x"FC90", x"FA10", x"F861", x"F72F", x"F66B", x"F6C6", x"F78E", x"F831", x"F918", x"F9FD", x"FA8B", x"FB1E", x"FBA2", x"FBAF", x"FBBF", x"FBCF", x"FB29", x"FA5F", x"F9AC", x"F85B", x"F70E", x"F69E", x"F5B4", x"F43E", x"F488", x"F61B", x"F7AB", x"FA14", x"FC88", x"FC89", x"FBED", x"FDDC", x"0125", x"04A8", x"097F", x"0DE0", x"0F9C", x"10DA", x"1273", x"120F", x"0FE2", x"0DC2", x"0AC4", x"072C", x"0518", x"03CD", x"01D1", x"0035", x"FEFD", x"FD06", x"FB8B", x"FB38", x"FAE1", x"FAC5", x"FBAE", x"FC4C", x"FC8D", x"FD86", x"FE54", x"FE34", x"FE6C", x"FE70", x"FD8D", x"FD25", x"FD66", x"FCE8", x"FC68", x"FC52", x"FAB5", x"F8AB", x"F875", x"F910", x"F951", x"FA48", x"F9F7", x"F695", x"F36C", x"F2D7", x"F35A", x"F52E", x"F8F5", x"FBED", x"FCFD", x"FEC6", x"009F", x"00D0", x"00A7", x"00BD", x"FFC7", x"FED3", x"FF00", x"FEC6", x"FDD8", x"FD3A", x"FC7E", x"FB85", x"FBF2", x"FD6B", x"FEDB", x"0095", x"01E8", x"01A6", x"00B9", x"FFF6", x"FEEB", x"FE91", x"FF88", x"00A6", x"020A", x"0457", x"0671", x"0829", x"0AB3", x"0C9C", x"0CA2", x"0CA9", x"0D2A", x"0CF7", x"0D4C", x"0EAE", x"0E16", x"0BED", x"0BA6", x"0D4F", x"0FC2", x"146B", x"19C5", x"1C71", x"1D9C", x"1F31", x"1F74", x"1E13", x"1CDD", x"1AE2", x"1790", x"153D", x"1440", x"12CC", x"1146", x"1003", x"0D9F", x"0A93", x"087D", x"06D3", x"0544", x"04F4", x"0551", x"05C5", x"0705", x"08FF", x"0ADE", x"0D21", x"0FCF", x"120F", x"1428", x"1628", x"1707", x"1739", x"1775", x"1640", x"136F", x"10D7", x"0E45", x"0B12", x"08C1", x"06CC", x"0292", x"FDD4", x"FBAE", x"FBA3", x"FD1E", x"0152", x"05ED", x"082B", x"09D2", x"0C0F", x"0CD3", x"0C17", x"0B8E", x"0A65", x"083B", x"0732", x"06EC", x"05C4", x"043E", x"0354", x"0249", x"0199", x"01F4", x"0281", x"02AE", x"02EE", x"0322", x"0327", x"035C", x"038E", x"039F", x"0416", x"0461", x"0458", x"04A5", x"04DD", x"04A7", x"056C", x"0706", x"0774", x"076F", x"0883", x"0978", x"0A59", x"0CCB", x"0E97", x"0D5A", x"0C23", x"0D07", x"0E72", x"10F3", x"1588", x"18D0", x"1998", x"1AD3", x"1C2B", x"1B26", x"18F5", x"168E", x"1296", x"0EAD", x"0D06", x"0C37", x"0AE4", x"0A01", x"08A6", x"0622", x"0422", x"02E5", x"019B", x"00FA", x"011D", x"00B2", x"0074", x"0119", x"01AA", x"028D", x"0496", x"0644", x"073D", x"08C0", x"09E2", x"09CA", x"0A2A", x"0A51", x"0862", x"067C", x"064B", x"0622", x"068E", x"0863", x"0879", x"0598", x"03A4", x"036A", x"038D", x"0585", x"090F", x"0AAC", x"0AD9", x"0C39", x"0D61", x"0D77", x"0E25", x"0EF8", x"0ED7", x"0F84", x"117A", x"12F9", x"141A", x"1551", x"154C", x"14A4", x"1494", x"145B", x"13E8", x"13E8", x"1315", x"10EA", x"0EC3", x"0CAF", x"0A70", x"097C", x"09B1", x"0987", x"09E3", x"0B16", x"0BCC", x"0CC6", x"0EFD", x"1033", x"0FC7", x"0FD1", x"0FB1", x"0EDF", x"0F82", x"10C2", x"0F4B", x"0C76", x"0AC6", x"095A", x"08ED", x"0B55", x"0DD9", x"0DFF", x"0DC1", x"0DCB", x"0C80", x"0B3A", x"0AD1", x"0955", x"0711", x"05ED", x"04F6", x"035B", x"021B", x"006E", x"FD54", x"FA4E", x"F826", x"F632", x"F557", x"F5EF", x"F6C0", x"F7E3", x"F9F5", x"FC06", x"FDEE", x"0040", x"023D", x"0376", x"04FA", x"062B", x"068D", x"0789", x"08D6", x"08CF", x"0834", x"07DA", x"0676", x"04F9", x"0515", x"04D0", x"0266", x"0030", x"FF37", x"FEC3", x"0079", x"04DD", x"089E", x"0A8B", x"0C76", x"0DE9", x"0DCF", x"0D89", x"0D4F", x"0BCF", x"09ED", x"090E", x"084E", x"0738", x"0659", x"058A", x"0480", x"03F9", x"0423", x"0492", x"0539", x"05F4", x"066A", x"06A8", x"064F", x"0535", x"0403", x"02CD", x"015C", x"004C", x"FFB2", x"FE75", x"FD5A", x"FDB4", x"FE79", x"FEDB", x"FFE8", x"0145", x"01B3", x"02CB", x"0530", x"0631", x"054F", x"0509", x"05B0", x"06C0", x"09FD", x"0EBF", x"11BE", x"12F1", x"1442", x"14A6", x"1350", x"1183", x"0F1F", x"0B46", x"0781", x"0527", x"032D", x"0137", x"FFC4", x"FE56", x"FCC7", x"FBAC", x"FB30", x"FB0D", x"FB8A", x"FC84", x"FDBC", x"FF35", x"0074", x"0119", x"019D", x"01EB", x"018B", x"012E", x"010A", x"0029", x"FF47", x"FF32", x"FEA9", x"FD29", x"FC4B", x"FBC6", x"FAE6", x"FB01", x"FBC7", x"FA4E", x"F703", x"F466", x"F29C", x"F1DB", x"F3FF", x"F7A1", x"F9E9", x"FB72", x"FD2D", x"FD95", x"FCD8", x"FC63", x"FB9B", x"FA3A", x"F98F", x"F9A0", x"F947", x"F91E", x"F94D", x"F97E", x"FA13", x"FB79", x"FCCB", x"FDFF", x"FF28", x"FF3F", x"FE87", x"FDD8", x"FD16", x"FC71", x"FCF1", x"FE33", x"FF6B", x"0174", x"0425", x"0694", x"0971", x"0CD8", x"0F11", x"1009", x"10C2", x"1080", x"0F6F", x"0F32", x"0EE6", x"0CD1", x"0A8E", x"096B", x"08DC", x"09EC", x"0D65", x"10B9", x"1261", x"139C", x"1441", x"1361", x"1249", x"112E", x"0EBF", x"0BB5", x"0946", x"0707", x"04E8", x"03D8", x"02DF", x"015E", x"FFF4", x"FEA1", x"FCE0", x"FB87", x"FAEB", x"FA72", x"FAB0", x"FC0C", x"FDD0", x"FFCE", x"024D", x"04C1", x"0723", x"09CB", x"0BD5", x"0CD8", x"0D33", x"0C85", x"0A66", x"0813", x"05B0", x"02AD", x"004F", x"FF2F", x"FD69", x"FA91", x"F86A", x"F6D4", x"F602", x"F7EF", x"FBF4", x"FEFD", x"00DF", x"0294", x"0332", x"02E1", x"0363", x"03B5", x"0284", x"00F6", x"FFD4", x"FE0E", x"FC42", x"FB41", x"FA16", x"F8A5", x"F7F5", x"F7D2", x"F75F", x"F71F", x"F714", x"F6D1", x"F6C5", x"F758", x"F7FA", x"F879", x"F916", x"F9A2", x"FA8F", x"FBC4", x"FCDE", x"FDF0", x"FF5D", x"0064", x"00E6", x"018C", x"01CA", x"0155", x"01D8", x"0337", x"035D", x"0273", x"01EC", x"014B", x"0127", x"036F", x"06C1", x"0851", x"08DA", x"096B", x"08C9", x"0756", x"0689", x"0525", x"023D", x"FF94", x"FDA9", x"FB0C", x"F826", x"F592", x"F278", x"EF2E", x"ECC9", x"EB29", x"E999", x"E8A4", x"E85D", x"E888", x"E972", x"EAEE", x"EC87", x"EE37", x"EFE1", x"F163", x"F326", x"F4BB", x"F566", x"F60F", x"F6CD", x"F6BB", x"F63F", x"F654", x"F5F4", x"F568", x"F663", x"F791", x"F68A", x"F484", x"F2C1", x"F095", x"EFCB", x"F20F", x"F4A4", x"F559", x"F5DD", x"F629", x"F536", x"F4E8", x"F60E", x"F6A5", x"F6C7", x"F7F8", x"F919", x"F971", x"FA57", x"FB48", x"FB54", x"FBA6", x"FC4B", x"FC28", x"FBB6", x"FB76", x"FA5C", x"F918", x"F884", x"F7CE", x"F700", x"F6FA", x"F70D", x"F6CF", x"F798", x"F8EC", x"FA16", x"FC3B", x"FF13", x"00FB", x"0297", x"0488", x"0574", x"05EA", x"073D", x"0751", x"04DA", x"0205", x"FF63", x"FCC4", x"FC71", x"FEB0", x"0027", x"0062", x"00D6", x"00B2", x"0005", x"00CB", x"01E1", x"0150", x"FFF7", x"FE48", x"FB4D", x"F82E", x"F616", x"F3ED", x"F1B8", x"F04B", x"EEAA", x"EC9B", x"EB2B", x"EA16", x"E90E", x"E90B", x"E9EE", x"EAA6", x"EBD1", x"ED40", x"EE24", x"EF2C", x"F0D0", x"F1DB", x"F2D5", x"F471", x"F56D", x"F57E", x"F609", x"F5F7", x"F4D8", x"F4EF", x"F5F8", x"F576", x"F3FF", x"F2A8", x"F012", x"EDF9", x"EF5B", x"F260", x"F476", x"F6BE", x"F8B0", x"F8CD", x"F91E", x"FAFE", x"FBB5", x"FADA", x"F9D3", x"F7DD", x"F4BE", x"F2C5", x"F1EE", x"F0CB", x"F061", x"F114", x"F177", x"F1B8", x"F25F", x"F20F", x"F09D", x"EF1F", x"ED2D", x"EAE0", x"E949", x"E83C", x"E77A", x"E7DC", x"E904", x"EA00", x"EBDF", x"EE86", x"F094", x"F278", x"F470", x"F4DB", x"F46A", x"F57E", x"F702", x"F78B", x"F864", x"F95A", x"F939", x"FA62", x"FE5D", x"0260", x"04F4", x"0729", x"080D", x"0735", x"070E", x"07E4", x"0788", x"0623", x"047E", x"01B6", x"FDF8", x"FADD", x"F81D", x"F581", x"F3D0", x"F2FF", x"F272", x"F263", x"F2B8", x"F34D", x"F44D", x"F560", x"F5A2", x"F57E", x"F4F9", x"F3E9", x"F381", x"F44E", x"F4A6", x"F4A9", x"F553", x"F57C", x"F498", x"F473", x"F43F", x"F29C", x"F1BA", x"F2DD", x"F370", x"F2F5", x"F2B5", x"F13D", x"EEA7", x"EEB7", x"F172", x"F393", x"F4E0", x"F592", x"F3E6", x"F124", x"F04F", x"F0C9", x"F101", x"F213", x"F34B", x"F34F", x"F329", x"F3D5", x"F477", x"F581", x"F783", x"F93F", x"FA35", x"FAD8", x"FAAA", x"F9BD", x"F92E", x"F896", x"F77D", x"F6EE", x"F6A6", x"F62A", x"F690", x"F7FD", x"F8E5", x"FA2F", x"FCB0", x"FEE9", x"00AF", x"0308", x"046A", x"03F1", x"03FF", x"04D8", x"048B", x"03F3", x"0410", x"0358", x"030F", x"05AE", x"09C3", x"0CC5", x"0F3B", x"107C", x"0F85", x"0E13", x"0DB3", x"0D05", x"0B9B", x"0A40", x"0831", x"0563", x"030F", x"0163", x"000E", x"FF81", x"FF39", x"FE51", x"FD1C", x"FB9B", x"F9C8", x"F8CE", x"F8F5", x"F93A", x"FA18", x"FBC9", x"FD35", x"FEB4", x"011B", x"02CA", x"02F4", x"0305", x"02BA", x"0129", x"000E", x"FFB6", x"FE0A", x"FC1C", x"FBE1", x"FBDA", x"FB26", x"FB11", x"FA5F", x"F7CF", x"F61A", x"F6DD", x"F816", x"F980", x"FB9C", x"FC90", x"FC59", x"FD3C", x"FF19", x"0068", x"016C", x"01E0", x"007F", x"FE38", x"FC48", x"FA89", x"F976", x"F99F", x"FA18", x"FA3B", x"FA50", x"F9CB", x"F8A9", x"F7FC", x"F790", x"F6F2", x"F6D7", x"F736", x"F74D", x"F7FA", x"F989", x"FA97", x"FB4D", x"FCA2", x"FD89", x"FDE6", x"FEF3", x"0002", x"FFED", x"0055", x"021A", x"03B3", x"0510", x"06B3", x"06E7", x"05C0", x"05D0", x"0797", x"0994", x"0BD1", x"0DE4", x"0E55", x"0DBF", x"0DD4", x"0E4D", x"0E41", x"0DE1", x"0C8F", x"0986", x"055D", x"00E4", x"FCAE", x"F994", x"F829", x"F810", x"F8F1", x"FA19", x"FB12", x"FC43", x"FDDC", x"FF56", x"00A1", x"01CB", x"020D", x"01AC", x"01F6", x"028B", x"02CE", x"0375", x"0445", x"040C", x"0381", x"0373", x"028C", x"00C2", x"FFFC", x"FFD4", x"FF37", x"FEF6", x"FEC4", x"FCF8", x"FAF5", x"FB12", x"FC9C", x"FE8D", x"0103", x"02BB", x"0266", x"01BA", x"0229", x"0301", x"0419", x"05C1", x"06B4", x"0675", x"05A7", x"0499", x"0350", x"02BD", x"0318", x"03D7", x"04C5", x"055E", x"0528", x"0495", x"03F1", x"02F4", x"020B", x"0177", x"00AE", x"0016", x"0088", x"0137", x"01DE", x"0353", x"0541", x"06DE", x"0905", x"0BA0", x"0CD1", x"0CE7", x"0D0F", x"0C8F", x"0B0A", x"09EE", x"08AC", x"066D", x"051B", x"061E", x"0803", x"0A0A", x"0C46", x"0D3B", x"0C92", x"0C10", x"0C4D", x"0C27", x"0B99", x"0A9B", x"0885", x"0575", x"025C", x"FF77", x"FD27", x"FBAF", x"FB08", x"FAA4", x"FA05", x"F897", x"F6D4", x"F57D", x"F49D", x"F458", x"F50D", x"F5F5", x"F671", x"F758", x"F8B0", x"F97D", x"FA62", x"FBD6", x"FCE3", x"FD93", x"FEFD", x"FFFF", x"FFB6", x"FF5B", x"FF74", x"FF0D", x"FE99", x"FE97", x"FD5D", x"FB05", x"F9DC", x"FA7F", x"FC43", x"FF5B", x"02E8", x"0529", x"0625", x"072A", x"0816", x"08B1", x"0943", x"0969", x"088E", x"06E5", x"04E5", x"0300", x"0211", x"0274", x"03E2", x"05C9", x"0705", x"06BA", x"0556", x"0378", x"0146", x"FF90", x"FED4", x"FE95", x"FE9B", x"FF88", x"00EA", x"0222", x"03D5", x"05F5", x"079A", x"08F4", x"0A38", x"0A82", x"09AA", x"0924", x"0920", x"0958", x"0A2D", x"0B6A", x"0B80", x"0AE3", x"0B0B", x"0C0C", x"0D7F", x"0F90", x"1186", x"123C", x"1250", x"12CC", x"136A", x"13DE", x"1449", x"1428", x"12BB", x"103A", x"0D26", x"09CD", x"0719", x"05B6", x"05C1", x"067F", x"0746", x"077A", x"0703", x"0620", x"050F", x"041D", x"0370", x"02A3", x"01F5", x"0190", x"0160", x"0153", x"01A6", x"01D5", x"0179", x"00EF", x"0078", x"FF95", x"FEE0", x"FF01", x"FF49", x"FF94", x"0023", x"0023", x"FE97", x"FCC2", x"FBB2", x"FAEF", x"FAA7", x"FAF0", x"FA75", x"F8B0", x"F758", x"F72A", x"F7B2", x"F949", x"FBB9", x"FD88", x"FE5B", x"FEBE", x"FE94", x"FE01", x"FE1D", x"FF20", x"0098", x"0259", x"03D9", x"0454", x"0403", x"0356", x"025A", x"01AB", x"015B", x"0114", x"00E6", x"0136", x"01A8", x"02B0", x"04D5", x"078A", x"0A60", x"0DCD", x"10D2", x"1271", x"135D", x"1421", x"1419", x"1421", x"1507", x"1526", x"1404", x"136E", x"13BA", x"1443", x"15BA", x"17C4", x"181E", x"170B", x"1651", x"15F5", x"158E", x"15EE", x"1670", x"15C5", x"1448", x"1290", x"106A", x"0E69", x"0D92", x"0DD9", x"0EE7", x"1021", x"10A8", x"1038", x"0F39", x"0DF8", x"0D2C", x"0D51", x"0DB3", x"0E02", x"0E82", x"0EBD", x"0E44", x"0E28", x"0E7F", x"0EAC", x"0F61", x"1102", x"120A", x"1217", x"1245", x"1231", x"119A", x"11DF", x"1281", x"1156", x"0ECE", x"0C73", x"0A4B", x"090B", x"09DA", x"0B89", x"0C19", x"0C1B", x"0C03", x"0B70", x"0ADA", x"0ACA", x"0A86", x"0988", x"07EF", x"05C4", x"0351", x"01A6", x"012E", x"0225", x"042A", x"05F4", x"06D6", x"0735", x"0738", x"06DC", x"06FF", x"0799", x"07BC", x"07B0", x"0808", x"0804", x"0792", x"07A9", x"07E1", x"07D2", x"0880", x"09E9", x"0ACC", x"0B7F", x"0C8D", x"0D43", x"0DC0", x"0F1D", x"1048", x"1036", x"0FC1", x"0FC5", x"0FE7", x"10E9", x"1315", x"14CD", x"1533", x"14F1", x"1444", x"1302", x"11D7", x"10AB", x"0EB4", x"0B9D", x"07A0", x"02DD", x"FE4F", x"FB38", x"FA05", x"FADE", x"FD10", x"FF43", x"00A6", x"0172", x"0187", x"0102", x"00A9", x"004D", x"FF81", x"FEA3", x"FE0A", x"FD54", x"FD0B", x"FD7C", x"FE23", x"FE9F", x"FF70", x"000B", x"0023", x"007B", x"011D", x"016D", x"021D", x"0375", x"0409", x"03A8", x"0343", x"02CF", x"0279", x"0386", x"0580", x"068A", x"067D", x"05FF", x"04B8", x"0360", x"0311", x"0356", x"033D", x"02F1", x"0241", x"00C9", x"FF7C", x"FF2C", x"FFD0", x"017A", x"03CC", x"0582", x"0621", x"05DC", x"04BA", x"035D", x"02AD", x"0287", x"0291", x"02D1", x"02F0", x"029D", x"02C6", x"03C2", x"051A", x"0747", x"0A3D", x"0C82", x"0DBF", x"0E86", x"0E1E", x"0CD0", x"0C8C", x"0D4B", x"0D65", x"0D41", x"0D60", x"0CF6", x"0CD4", x"0E8A", x"10A3", x"113C", x"1108", x"105C", x"0EE0", x"0DA5", x"0D85", x"0D40", x"0C15", x"0A6C", x"07FC", x"0494", x"012E", x"FE56", x"FC54", x"FB3D", x"FAA2", x"F9C8", x"F88F", x"F6FD", x"F553", x"F47C", x"F49A", x"F500", x"F5C4", x"F70B", x"F7E6", x"F8BC", x"FA50", x"FBD2", x"FCF6", x"FEAB", x"008E", x"0135", x"0136", x"00E3", x"FF39", x"FD40", x"FCC8", x"FCB8", x"FB9F", x"FA72", x"F971", x"F859", x"F8C9", x"FBCA", x"FF2D", x"016F", x"032F", x"0445", x"0488", x"0516", x"063A", x"06D1", x"066C", x"0537", x"02FD", x"0004", x"FD29", x"FB28", x"FA52", x"FA3B", x"F9DC", x"F8C8", x"F733", x"F516", x"F336", x"F26C", x"F22B", x"F1AF", x"F1A0", x"F1DD", x"F1D4", x"F219", x"F32A", x"F404", x"F4B0", x"F62C", x"F7B2", x"F85E", x"F8F3", x"F959", x"F8E6", x"F8AE", x"F9C1", x"FA8B", x"FA61", x"FA2B", x"F9EC", x"F99C", x"FAD6", x"FD91", x"FFCC", x"00FB", x"01A4", x"019F", x"013B", x"019E", x"0293", x"0333", x"0334", x"022C", x"FFBD", x"FC84", x"F983", x"F77E", x"F71C", x"F7F2", x"F8BB", x"F918", x"F8FA", x"F800", x"F6BA", x"F5FA", x"F55F", x"F487", x"F424", x"F3F1", x"F318", x"F263", x"F235", x"F1E8", x"F1FC", x"F303", x"F3EC", x"F423", x"F470", x"F45D", x"F39E", x"F3A4", x"F47E", x"F47E", x"F387", x"F22E", x"EFC3", x"ED1A", x"EC2A", x"EC55", x"EC12", x"EBD5", x"EBBE", x"EB1C", x"EAEC", x"EC44", x"EDF5", x"EF69", x"F0E4", x"F1B8", x"F160", x"F0F6", x"F0E7", x"F123", x"F248", x"F430", x"F5AF", x"F680", x"F6A3", x"F58B", x"F3B1", x"F211", x"F0B3", x"EF92", x"EF2E", x"EF0A", x"EED3", x"EF66", x"F0E3", x"F309", x"F65A", x"FA76", x"FE09", x"00F2", x"035E", x"044F", x"0465", x"0539", x"0611", x"05CF", x"0522", x"03D9", x"0156", x"FF7C", x"FFD3", x"008F", x"00AD", x"00CF", x"006B", x"FF47", x"FF2D", x"006E", x"0164", x"01CB", x"0201", x"014B", x"FFE0", x"FEEF", x"FE99", x"FEA7", x"FF70", x"006D", x"00B3", x"0041", x"FF05", x"FD02", x"FB0D", x"F960", x"F7A5", x"F638", x"F525", x"F3E8", x"F31E", x"F370", x"F411", x"F50C", x"F71D", x"F951", x"FA93", x"FBBB", x"FC65", x"FB8B", x"FACA", x"FB8B", x"FC07", x"FB42", x"FA39", x"F827", x"F512", x"F3ED", x"F582", x"F71D", x"F7FC", x"F8B3", x"F833", x"F6BD", x"F687", x"F768", x"F782", x"F759", x"F740", x"F623", x"F46A", x"F338", x"F279", x"F236", x"F324", x"F4B0", x"F5F4", x"F6D1", x"F705", x"F66F", x"F5CA", x"F529", x"F453", x"F3B1", x"F35A", x"F2B2", x"F262", x"F2BD", x"F325", x"F3EE", x"F5EC", x"F82D", x"F9DC", x"FBBC", x"FD19", x"FD49", x"FDEA", x"FFCB", x"00F5", x"012F", x"014C", x"006C", x"FF12", x"FFBE", x"0217", x"03CF", x"04F6", x"05B8", x"04E2", x"0324", x"0218", x"00EC", x"FEE9", x"FD06", x"FB05", x"F83B", x"F575", x"F35E", x"F1DA", x"F1AC", x"F308", x"F4D7", x"F6B8", x"F883", x"F93B", x"F926", x"F902", x"F86F", x"F78B", x"F76E", x"F78F", x"F707", x"F69E", x"F63A", x"F4F7", x"F428", x"F496", x"F4CD", x"F4BF", x"F51F", x"F4A8", x"F361", x"F396", x"F4DF", x"F564", x"F5DB", x"F65E", x"F59A", x"F54E", x"F7AA", x"FABA", x"FCCF", x"FEB8", x"FF74", x"FE2E", x"FD3B", x"FD87", x"FD43", x"FCB1", x"FCA7", x"FBDB", x"FA43", x"F98C", x"F910", x"F836", x"F832", x"F8F0", x"F93C", x"F9C8", x"FA9A", x"FA5D", x"F973", x"F8E1", x"F80F", x"F733", x"F729", x"F71C", x"F68E", x"F692", x"F72D", x"F80E", x"FA08", x"FCA6", x"FE6F", x"FFA6", x"0076", x"FFFC", x"FF6A", x"0049", x"015B", x"01C3", x"0220", x"0174", x"FF3E", x"FE32", x"FF42", x"008A", x"01AD", x"02F5", x"029E", x"00FA", x"0059", x"006A", x"FFD2", x"FF54", x"FEBB", x"FCC3", x"FA43", x"F847", x"F634", x"F433", x"F340", x"F2A4", x"F1D0", x"F141", x"F08E", x"EF45", x"EE3B", x"ED82", x"ECD2", x"ECA7", x"ECFC", x"ED25", x"EDAF", x"EED0", x"EFAD", x"F0C6", x"F2AC", x"F46A", x"F580", x"F6DA", x"F729", x"F5D1", x"F4FC", x"F597", x"F5D9", x"F624", x"F6B2", x"F582", x"F345", x"F369", x"F5B6", x"F820", x"FB16", x"FDF8", x"FE8F", x"FE36", x"FF29", x"000E", x"0019", x"00AD", x"0143", x"0089", x"FFAB", x"FEEC", x"FCE1", x"FA32", x"F858", x"F6F1", x"F60A", x"F64E", x"F6BB", x"F67A", x"F608", x"F594", x"F4C7", x"F47B", x"F4CC", x"F535", x"F639", x"F7EF", x"F9B7", x"FBD5", x"FEA4", x"00F5", x"02B1", x"0449", x"04B5", x"03C9", x"0357", x"035A", x"027A", x"0150", x"000D", x"FD55", x"FA9F", x"FA44", x"FB4E", x"FC4C", x"FE0C", x"FFA9", x"FFED", x"004D", x"01E0", x"0316", x"03D2", x"0504", x"059A", x"04F6", x"0406", x"02B6", x"0094", x"FEF3", x"FE4D", x"FE14", x"FE40", x"FEB0", x"FE50", x"FD4B", x"FC3C", x"FACA", x"F967", x"F8BE", x"F82C", x"F781", x"F76B", x"F749", x"F6BA", x"F6F5", x"F7CC", x"F83B", x"F8DB", x"F9B1", x"F918", x"F7FE", x"F832", x"F873", x"F7D1", x"F72D", x"F556", x"F165", x"EE57", x"EDF3", x"EE64", x"EF63", x"F135", x"F1A0", x"F051", x"F010", x"F0C7", x"F121", x"F230", x"F400", x"F4D4", x"F53B", x"F66B", x"F6EE", x"F6A1", x"F70B", x"F7B9", x"F83F", x"F9A9", x"FB7C", x"FC30", x"FC3F", x"FC48", x"FBB5", x"FB2B", x"FB6D", x"FB74", x"FB32", x"FB8E", x"FC81", x"FE14", x"012F", x"0504", x"0868", x"0B93", x"0DFA", x"0ECD", x"0F75", x"10CE", x"11CE", x"124C", x"12A1", x"1143", x"0E5E", x"0C6C", x"0BE5", x"0BA8", x"0C44", x"0D4B", x"0CF0", x"0BC4", x"0B53", x"0ABB", x"097A", x"08A5", x"07F4", x"068F", x"05AD", x"0591", x"0554", x"0547", x"061F", x"073F", x"0867", x"09FF", x"0B2F", x"0B4F", x"0AEE", x"0A0A", x"08B8", x"078A", x"0692", x"05A4", x"052C", x"052B", x"051D", x"0578", x"0646", x"06DA", x"07AF", x"0927", x"09F6", x"09FC", x"0AB5", x"0BD2", x"0C7F", x"0D77", x"0E03", x"0C3E", x"0982", x"0854", x"0826", x"0888", x"0A40", x"0BA9", x"0AE2", x"0999", x"08DB", x"0756", x"0585", x"04C2", x"0422", x"034A", x"03C1", x"04DE", x"0506", x"04F6", x"0569", x"0593", x"062F", x"07F9", x"0990", x"0A24", x"0A64", x"0A17", x"0915", x"0828", x"0777", x"066C", x"0592", x"057A", x"05CB", x"06E9", x"08DE", x"0AAF", x"0C52", x"0DE6", x"0EB0", x"0EE5", x"0FDF", x"1120", x"11C3", x"122B", x"11BE", x"0F60", x"0CF0", x"0C4F", x"0C9F", x"0D72", x"0F1F", x"0FFE", x"0EDD", x"0D73", x"0C3A", x"0A2A", x"081E", x"0717", x"05DF", x"047B", x"03D0", x"0313", x"01C2", x"011E", x"0175", x"022B", x"036D", x"0502", x"0576", x"04E6", x"0412", x"02F4", x"0205", x"01D6", x"01AB", x"0150", x"0110", x"00A7", x"001A", x"001D", x"0056", x"0041", x"0081", x"00BD", x"0002", x"FF8C", x"004C", x"0138", x"0251", x"03ED", x"0429", x"02A7", x"01F1", x"02D4", x"0444", x"06F7", x"0A4E", x"0BB0", x"0B48", x"0AFF", x"0A0F", x"083C", x"0727", x"065A", x"04C5", x"03C2", x"03B1", x"02E4", x"0190", x"009D", x"FF29", x"FD9F", x"FD9C", x"FE7A", x"FF0D", x"000A", x"012E", x"01AB", x"026C", x"03E5", x"04F0", x"059E", x"06B1", x"07A4", x"08B7", x"0ACA", x"0D1F", x"0F0B", x"1104", x"1264", x"129D", x"12DF", x"1391", x"13DF", x"1417", x"1464", x"1342", x"1146", x"1074", x"10B3", x"116D", x"134B", x"154C", x"15B5", x"1573", x"156D", x"148D", x"12F4", x"118E", x"0F84", x"0CB3", x"0A68", x"088E", x"063D", x"03FE", x"0232", x"0007", x"FE38", x"FD5D", x"FCC3", x"FBF9", x"FBA2", x"FB68", x"FB18", x"FB46", x"FBBB", x"FBE1", x"FC00", x"FC5A", x"FCA5", x"FD5E", x"FE6C", x"FF46", x"0003", x"00CC", x"00B4", x"0030", x"002B", x"006F", x"00D4", x"01EF", x"028E", x"0145", x"FF6A", x"FE81", x"FE3B", x"FF6B", x"0280", x"054D", x"068E", x"077C", x"07FC", x"076B", x"070F", x"0784", x"075B", x"0722", x"07AE", x"07D9", x"06D9", x"05E2", x"0476", x"0238", x"00B9", x"0052", x"FFC5", x"FF27", x"FEF5", x"FE1B", x"FCEA", x"FC71", x"FC0E", x"FB2D", x"FABB", x"FAC9", x"FB19", x"FCB9", x"FF9B", x"0296", x"0584", x"084D", x"09C1", x"0A7F", x"0BBF", x"0CE5", x"0DA2", x"0E50", x"0DA9", x"0AB1", x"078E", x"058A", x"044D", x"04B4", x"06EB", x"089C", x"0943", x"0A13", x"0A72", x"09C9", x"097B", x"097D", x"08AC", x"0807", x"0832", x"07D2", x"0732", x"071B", x"06BF", x"0605", x"060F", x"0641", x"0591", x"049B", x"0357", x"0108", x"FECD", x"FD3B", x"FB89", x"F9FB", x"F940", x"F8BA", x"F8B1", x"F9BB", x"FB18", x"FC29", x"FD82", x"FE6F", x"FE6E", x"FEAA", x"FF65", x"FFB1", x"0022", x"0086", x"FEF7", x"FBE0", x"F932", x"F6FD", x"F58E", x"F649", x"F7EB", x"F867", x"F8A1", x"F91B", x"F8CB", x"F8AD", x"F9AA", x"FA39", x"FA2B", x"FAEE", x"FBDC", x"FC41", x"FD43", x"FE3D", x"FDC3", x"FD13", x"FD0D", x"FCC6", x"FC92", x"FD2E", x"FD0A", x"FBD2", x"FB05", x"FA61", x"F961", x"F960", x"FA6C", x"FBC2", x"FE3D", x"0245", x"064A", x"0A27", x"0E10", x"1086", x"11AD", x"12DC", x"13F3", x"1472", x"154E", x"158A", x"135C", x"1014", x"0D03", x"0A13", x"085E", x"08CE", x"0989", x"0954", x"092E", x"08B6", x"0748", x"0648", x"05CF", x"04BE", x"03B1", x"0399", x"0395", x"03C7", x"050D", x"0651", x"0703", x"0803", x"0911", x"0946", x"0942", x"092E", x"0833", x"06F5", x"064F", x"056C", x"0436", x"032D", x"0200", x"00A5", x"003B", x"0084", x"0102", x"021A", x"0365", x"03D6", x"042E", x"04E9", x"0593", x"06BF", x"08DB", x"0A09", x"095F", x"080C", x"063E", x"0467", x"044D", x"05EB", x"072B", x"07AC", x"07B5", x"063B", x"03CA", x"021A", x"00C5", x"FF65", x"FF0F", x"FF7E", x"FFA4", x"003A", x"014B", x"0175", x"0102", x"0112", x"00F6", x"00D5", x"01CB", x"02FC", x"035E", x"03BA", x"0415", x"0361", x"026A", x"01DC", x"00FE", x"0072", x"014B", x"02B3", x"0427", x"0637", x"07F2", x"0890", x"098B", x"0B3E", x"0CF3", x"0F49", x"11E9", x"1299", x"1141", x"0F96", x"0DC6", x"0C66", x"0D26", x"0F0E", x"1029", x"10D7", x"1129", x"100C", x"0E36", x"0CC3", x"0AAE", x"0831", x"06A1", x"05AD", x"0518", x"05FC", x"07B0", x"08CB", x"09AF", x"0A72", x"0A1C", x"095D", x"092D", x"088A", x"0781", x"071E", x"06BB", x"05B1", x"04D6", x"03F4", x"0272", x"015B", x"0111", x"008B", x"0015", x"FFEE", x"FF21", x"FE1F", x"FE3A", x"FEF4", x"0015", x"023C", x"03F4", x"0390", x"01F5", x"FFE8", x"FD84", x"FC7D", x"FDDF", x"FFE5", x"017F", x"02F6", x"030B", x"0197", x"0041", x"FF22", x"FD8D", x"FC55", x"FB9B", x"FA38", x"F8EE", x"F86D", x"F763", x"F59E", x"F45F", x"F319", x"F1E8", x"F240", x"F3BE", x"F4C0", x"F5B2", x"F6D1", x"F6F4", x"F6A5", x"F6E0", x"F6DE", x"F6E1", x"F831", x"FA7B", x"FD02", x"0040", x"0356", x"04EC", x"05CB", x"0686", x"06B3", x"0748", x"08E1", x"09AF", x"08E6", x"074B", x"04FD", x"0275", x"01C9", x"0336", x"050D", x"0702", x"08DB", x"095E", x"08D1", x"0850", x"0758", x"05AE", x"041D", x"0266", x"0020", x"FE43", x"FCE4", x"FB33", x"F96E", x"F7F0", x"F613", x"F409", x"F2C1", x"F1B6", x"F09F", x"F035", x"F047", x"F01E", x"EFF4", x"EFC0", x"EF28", x"EEB6", x"EF04", x"EF99", x"F063", x"F165", x"F1F9", x"F208", x"F23B", x"F27A", x"F2A2", x"F37D", x"F499", x"F4B5", x"F3C9", x"F27D", x"F0E3", x"F02D", x"F1C2", x"F4F5", x"F86A", x"FBBD", x"FE1F", x"FEE4", x"FEC0", x"FE86", x"FE1A", x"FDE6", x"FE3A", x"FE8A", x"FE94", x"FEC7", x"FEA4", x"FDB4", x"FC47", x"FA4E", x"F78C", x"F535", x"F40E", x"F3D2", x"F467", x"F5DA", x"F6F5", x"F706", x"F678", x"F56B", x"F42C", x"F3E9", x"F533", x"F748", x"F9FD", x"FCD5", x"FEA2", x"FF5A", x"FFDA", x"0013", x"0049", x"0115", x"01A1", x"0057", x"FD87", x"FA07", x"F647", x"F3BA", x"F3B2", x"F53F", x"F73D", x"F99B", x"FBC5", x"FCCF", x"FD2F", x"FD24", x"FC6C", x"FB71", x"FAE0", x"FA79", x"FA67", x"FB10", x"FBF7", x"FCD1", x"FD6F", x"FD66", x"FC10", x"FA3F", x"F82F", x"F5A0", x"F343", x"F199", x"F030", x"EEFE", x"EE5D", x"EDDC", x"ED47", x"ED5A", x"EE26", x"EF0A", x"F008", x"F0B6", x"F07E", x"EFE4", x"EFBE", x"F028", x"F160", x"F363", x"F4D1", x"F45E", x"F255", x"EF09", x"EB47", x"E8AD", x"E826", x"E903", x"EAB2", x"ECC7", x"EE36", x"EE86", x"EE17", x"ED39", x"EC60", x"EC2A", x"ECA8", x"ED6F", x"EEA3", x"EFCA", x"F073", x"F0AC", x"F068", x"EF4D", x"EDF6", x"ED60", x"ED25", x"ED0C", x"ED39", x"ED2C", x"EC5A", x"EB50", x"EA79", x"E9C0", x"E9BF", x"EB38", x"EDC4", x"F0FB", x"F46F", x"F747", x"F907", x"FA4C", x"FB6F", x"FCB0", x"FEB3", x"0124", x"02B6", x"02D2", x"0184", x"FEE8", x"FC0B", x"FA6E", x"FA4A", x"FAD3", x"FBA4", x"FC4C", x"FC22", x"FB72", x"FAB7", x"FA1B", x"F98F", x"F93C", x"F8F0", x"F888", x"F879", x"F8DE", x"F9E5", x"FB69", x"FD1D", x"FE40", x"FEF4", x"FF5A", x"FF61", x"FF41", x"FF3A", x"FF30", x"FEB6", x"FDB4", x"FC42", x"FA78", x"F8EC", x"F82D", x"F846", x"F8AF", x"F90E", x"F91E", x"F922", x"F97C", x"FA6F", x"FC25", x"FE74", x"008D", x"016A", x"009D", x"FE58", x"FB19", x"F848", x"F70A", x"F762", x"F85E", x"F96D", x"F9F3", x"F95F", x"F7AE", x"F5AF", x"F3D2", x"F265", x"F1EC", x"F27F", x"F390", x"F4B9", x"F601", x"F73A", x"F823", x"F86B", x"F834", x"F788", x"F6E7", x"F6E9", x"F7C3", x"F945", x"FAAC", x"FB4E", x"FAC1", x"F917", x"F709", x"F575", x"F4F8", x"F595", x"F724", x"F8FB", x"FAC8", x"FC88", x"FE5A", x"0017", x"022E", x"04A8", x"06D9", x"07C8", x"0776", x"05ED", x"0388", x"01BA", x"017B", x"0244", x"0358", x"0492", x"055B", x"04D2", x"0327", x"00C2", x"FDD7", x"FAEB", x"F912", x"F86B", x"F8A3", x"F97C", x"FB13", x"FCEF", x"FEA6", x"FFAE", x"FFDB", x"FF27", x"FDD7", x"FC85", x"FBAE", x"FB41", x"FAF4", x"FABF", x"FA5E", x"F990", x"F885", x"F7AA", x"F6FB", x"F660", x"F5D3", x"F505", x"F3C6", x"F2B2", x"F249", x"F2BA", x"F48B", x"F753", x"F9CB", x"FAEC", x"FA65", x"F877", x"F5F3", x"F4A1", x"F547", x"F781", x"FA9B", x"FDEF", x"0071", x"0125", x"001E", x"FDC9", x"FAB9", x"F790", x"F502", x"F320", x"F174", x"EFC4", x"EE8E", x"EDB8", x"ECD0", x"EBCB", x"EB27", x"EAE9", x"EB6E", x"ED46", x"F030", x"F316", x"F595", x"F755", x"F816", x"F817", x"F855", x"F936", x"FAE5", x"FD55", x"FFD9", x"01BF", x"0321", x"0435", x"0519", x"0672", x"0876", x"0A86", x"0BE0", x"0C36", x"0AF8", x"0860", x"0600", x"04FB", x"05AA", x"07BA", x"0A58", x"0C35", x"0CAA", x"0BB2", x"09B8", x"0770", x"056F", x"03AC", x"0212", x"008B", x"FEBA", x"FCF9", x"FC0E", x"FBE1", x"FBE0", x"FBDE", x"FBB9", x"FB13", x"FA60", x"FA43", x"FA7A", x"FAD3", x"FB4E", x"FB60", x"FAD1", x"F9FD", x"F92C", x"F870", x"F81B", x"F800", x"F76C", x"F6C6", x"F699", x"F6BF", x"F750", x"F8DF", x"FAF1", x"FCC0", x"FE57", x"FF43", x"FEBC", x"FD41", x"FC5A", x"FC9A", x"FE3D", x"0118", x"043F", x"0678", x"0761", x"06FA", x"05AA", x"0417", x"02CA", x"0224", x"0260", x"02F0", x"033E", x"0379", x"03BD", x"0386", x"02EB", x"0223", x"00B6", x"FEE7", x"FDE0", x"FDD5", x"FE52", x"FF54", x"0035", x"FFC0", x"FE40", x"FCA8", x"FB28", x"FA23", x"FA92", x"FBB2", x"FCDE", x"FEC1", x"0163", x"03B2", x"05C4", x"0812", x"09CA", x"0A90", x"0AE6", x"0A13", x"0754", x"03B2", x"00C5", x"FF17", x"FF1A", x"00D0", x"033B", x"053F", x"067D", x"06B8", x"062A", x"053D", x"0451", x"03F2", x"0467", x"04F9", x"0583", x"0689", x"0805", x"0909", x"09BC", x"09A6", x"07CF", x"04C3", x"022A", x"0010", x"FE5C", x"FDB9", x"FD7E", x"FC9F", x"FBC1", x"FB8C", x"FB57", x"FB8D", x"FCAA", x"FDCE", x"FE69", x"FF4E", x"0052", x"00A3", x"014C", x"02DD", x"0472", x"05DC", x"06E1", x"060B", x"02E3", x"FF16", x"FC14", x"FAB5", x"FBA3", x"FE64", x"0166", x"03BF", x"04C6", x"0434", x"02CC", x"013E", x"FFE3", x"FF40", x"FF74", x"FF48", x"FEB5", x"FE9D", x"FE95", x"FE03", x"FD82", x"FCD2", x"FB21", x"F9C4", x"F9E1", x"FAA6", x"FBBF", x"FD7E", x"FEAD", x"FECF", x"FF21", x"000B", x"012E", x"0354", x"0675", x"0907", x"0B2D", x"0D7B", x"0F27", x"1035", x"11D9", x"13A9", x"14D9", x"160D", x"1690", x"14EE", x"11AF", x"0E57", x"0B82", x"0A33", x"0B6E", x"0DBF", x"0FC6", x"10FE", x"10DD", x"0F4E", x"0DD4", x"0D07", x"0C9E", x"0D03", x"0DBB", x"0DBC", x"0DAB", x"0E94", x"0FE6", x"1152", x"133D", x"146F", x"1453", x"1432", x"1459", x"1411", x"1406", x"1428", x"132C", x"1168", x"0FAA", x"0D5A", x"0AA5", x"08B6", x"06D0", x"0492", x"0393", x"043D", x"0562", x"0799", x"0AFA", x"0DB4", x"0FA5", x"11CF", x"12E8", x"11CC", x"0FC8", x"0DB7", x"0BC5", x"0B7C", x"0D41", x"0F43", x"104A", x"1016", x"0E11", x"0AB9", x"077F", x"0500", x"0386", x"038F", x"044C", x"050B", x"062C", x"078B", x"0893", x"09BF", x"0AE1", x"0AD1", x"0A11", x"09AE", x"095F", x"0972", x"0AA5", x"0BC0", x"0B6B", x"0A78", x"0909", x"06C2", x"051E", x"0512", x"053F", x"05D4", x"081A", x"0B22", x"0DE0", x"1144", x"14CB", x"1724", x"191F", x"1B5E", x"1C26", x"1AC4", x"1877", x"15C3", x"134B", x"127B", x"1361", x"146D", x"14C4", x"1409", x"11FE", x"0F18", x"0C2B", x"09B8", x"0891", x"0896", x"090D", x"09EB", x"0B74", x"0D06", x"0E97", x"106F", x"1135", x"0FBB", x"0D20", x"0A23", x"06E9", x"04E9", x"04D0", x"0507", x"04E5", x"050C", x"04CD", x"03D0", x"036F", x"03B2", x"037C", x"0381", x"04C9", x"061E", x"0757", x"0975", x"0BE4", x"0DE1", x"101B", x"1216", x"11B9", x"0EEB", x"0B22", x"0766", x"0510", x"057D", x"080E", x"0B0B", x"0D54", x"0E38", x"0D65", x"0B5A", x"08C8", x"0662", x"04E2", x"03F3", x"02EE", x"01EC", x"00E4", x"FF85", x"FE3D", x"FD86", x"FCB1", x"FB8A", x"FB37", x"FBCA", x"FCDF", x"FEE5", x"016A", x"0303", x"039A", x"03D5", x"036B", x"02E2", x"035D", x"049B", x"05E0", x"07D5", x"0A58", x"0C56", x"0E0E", x"1005", x"1176", x"127B", x"13B6", x"1469", x"135A", x"1117", x"0E93", x"0C6D", x"0BD4", x"0D7F", x"1050", x"12ED", x"1489", x"149D", x"131D", x"10E0", x"0EA7", x"0CFE", x"0C1B", x"0B75", x"0A79", x"095E", x"083A", x"0745", x"0711", x"077D", x"07BC", x"0794", x"0753", x"069D", x"05CD", x"058B", x"0578", x"0521", x"04C5", x"041C", x"028E", x"00D2", x"FF43", x"FD34", x"FB1B", x"FA12", x"F9DA", x"FA11", x"FB84", x"FD95", x"FF1C", x"00A3", x"02AF", x"03EE", x"03B2", x"02ED", x"01EB", x"012E", x"0254", x"05B8", x"09A5", x"0CC8", x"0EA1", x"0E8F", x"0CA5", x"0A1D", x"07ED", x"0660", x"05A0", x"0597", x"05C2", x"05B0", x"0550", x"04D3", x"044C", x"0392", x"0285", x"013F", x"FFA0", x"FE02", x"FD38", x"FD83", x"FE4E", x"FF12", x"FF4E", x"FE20", x"FBCC", x"F9C3", x"F86C", x"F7BE", x"F855", x"FA5E", x"FCC3", x"FF23", x"01D2", x"040C", x"054E", x"066F", x"07A0", x"0773", x"0578", x"02A0", x"FF81", x"FCD8", x"FC26", x"FDA8", x"FFA0", x"00FB", x"01B2", x"018C", x"002B", x"FE90", x"FD9C", x"FD34", x"FD4D", x"FE4A", x"FFAE", x"00AD", x"017B", x"02AB", x"03DE", x"0485", x"0493", x"0395", x"0124", x"FE2E", x"FBF7", x"FABD", x"FA1C", x"FA25", x"FA1F", x"F94B", x"F823", x"F779", x"F704", x"F675", x"F67E", x"F70E", x"F74D", x"F77A", x"F816", x"F8A1", x"F91F", x"FA85", x"FC5D", x"FCA4", x"FB07", x"F889", x"F59A", x"F39A", x"F44A", x"F751", x"FAB4", x"FD9D", x"FFEC", x"00A1", x"FFC2", x"FE68", x"FD08", x"FB96", x"FADD", x"FB02", x"FB5A", x"FB7F", x"FB91", x"FB74", x"FAFF", x"FA84", x"F9F2", x"F94A", x"F8AE", x"F86D", x"F8BC", x"F9B1", x"FB10", x"FC88", x"FDE0", x"FEDA", x"FF92", x"0089", x"01C0", x"0312", x"04F0", x"072F", x"0912", x"0A8C", x"0BE9", x"0CBA", x"0D1B", x"0DE1", x"0E49", x"0CFD", x"0A4E", x"0750", x"0475", x"02F7", x"040A", x"069E", x"08EB", x"0AB6", x"0BAA", x"0B16", x"09A1", x"088E", x"07F7", x"07E3", x"08AD", x"09BD", x"0A1E", x"09CF", x"0948", x"08A2", x"082A", x"081F", x"0831", x"07F5", x"077F", x"0717", x"06EE", x"0701", x"073B", x"0735", x"0648", x"0454", x"01F1", x"FF5B", x"FC92", x"FA4E", x"F937", x"F8CF", x"F90A", x"FA3E", x"FBA8", x"FC6D", x"FD87", x"FF17", x"FFDD", x"FF3F", x"FDE6", x"FB9D", x"F911", x"F882", x"FA4D", x"FCF6", x"FF7D", x"018F", x"01DF", x"0066", x"FE9D", x"FCFA", x"FB70", x"FA8F", x"FA92", x"FA87", x"FA59", x"FA55", x"FA50", x"FA26", x"FA38", x"FA45", x"F9DF", x"F8E6", x"F7CC", x"F6EF", x"F6D2", x"F7C7", x"F96B", x"FAF8", x"FB80", x"FB01", x"FA1D", x"F932", x"F8BC", x"F961", x"FB39", x"FD53", x"FF9D", x"020F", x"03D2", x"04A7", x"059D", x"068F", x"060E", x"040F", x"0119", x"FD4C", x"F9B5", x"F868", x"F94B", x"FAA5", x"FBCF", x"FC75", x"FB93", x"F921", x"F68C", x"F465", x"F2A5", x"F235", x"F372", x"F549", x"F6EF", x"F87F", x"F9C9", x"FA58", x"FA91", x"FA90", x"F9AD", x"F7B1", x"F597", x"F419", x"F331", x"F339", x"F3FE", x"F44B", x"F384", x"F277", x"F19C", x"F098", x"EFED", x"F057", x"F129", x"F210", x"F39A", x"F55F", x"F62C", x"F6B3", x"F804", x"F955", x"F9AF", x"F957", x"F7F9", x"F55F", x"F369", x"F3B3", x"F586", x"F7C8", x"FA3F", x"FBDE", x"FBC9", x"FA84", x"F8D3", x"F68D", x"F411", x"F22C", x"F0A9", x"EF25", x"EDAE", x"EC44", x"EAD9", x"E9AB", x"E90F", x"E8E7", x"E914", x"E987", x"EA41", x"EB63", x"ECD8", x"EE77", x"F009", x"F12B", x"F1AC", x"F217", x"F2C8", x"F3A7", x"F503", x"F728", x"F99F", x"FBD7", x"FE0D", x"FFCE", x"007D", x"00E0", x"01BD", x"021D", x"0146", x"FF7B", x"FCF3", x"F9EC", x"F870", x"F96F", x"FBD1", x"FE51", x"009C", x"0193", x"008B", x"FE43", x"FBD3", x"F96D", x"F7D5", x"F7B9", x"F88E", x"F944", x"F9AD", x"F9E8", x"F9E9", x"F9F6", x"FA61", x"FABC", x"FA4B", x"F94F", x"F83B", x"F733", x"F662", x"F602", x"F552", x"F372", x"F0CA", x"EE07", x"EB16", x"E87C", x"E719", x"E6B7", x"E6D9", x"E7EF", x"E9DE", x"EB45", x"EC36", x"EDB0", x"EF99", x"F139", x"F2CE", x"F3E7", x"F381", x"F2A0", x"F2D5", x"F42C", x"F5F1", x"F7E4", x"F924", x"F880", x"F657", x"F38E", x"F08C", x"EDFB", x"EC9F", x"EC78", x"ECCE", x"ED86", x"EE49", x"EEF0", x"EF91", x"F067", x"F12D", x"F1A8", x"F1BF", x"F168", x"F0E0", x"F08A", x"F0A6", x"F12B", x"F19D", x"F17A", x"F0C5", x"EFC4", x"EEAE", x"EDF2", x"EE0D", x"EED6", x"EFD3", x"F153", x"F317", x"F478", x"F5AA", x"F782", x"F981", x"FAA5", x"FADB", x"F9E6", x"F774", x"F4C6", x"F3A8", x"F409", x"F4FC", x"F675", x"F800", x"F85B", x"F788", x"F65D", x"F4B7", x"F2CC", x"F1E1", x"F277", x"F383", x"F4CB", x"F62B", x"F6FA", x"F6FA", x"F6FE", x"F6E3", x"F629", x"F4F1", x"F3C1", x"F285", x"F1A9", x"F1C9", x"F27A", x"F2B3", x"F276", x"F20E", x"F16E", x"F0C5", x"F0B1", x"F0FD", x"F113", x"F11E", x"F186", x"F1A9", x"F11D", x"F0B0", x"F0E9", x"F140", x"F18A", x"F1C8", x"F116", x"EF4C", x"EE1C", x"EEB4", x"F06B", x"F2F1", x"F5FE", x"F836", x"F8DA", x"F889", x"F785", x"F58B", x"F35B", x"F1D3", x"F097", x"EFB1", x"EF59", x"EF10", x"EEAE", x"EEA4", x"EF04", x"EFA8", x"F0E0", x"F277", x"F3F5", x"F57D", x"F741", x"F8F3", x"FA99", x"FC40", x"FD4F", x"FDDC", x"FE4D", x"FE97", x"FEE1", x"FFC2", x"00DF", x"01B8", x"02A4", x"0348", x"02F5", x"02C7", x"03B1", x"0489", x"04BD", x"049E", x"0343", x"00C4", x"FF9B", x"00BD", x"02C9", x"0571", x"0899", x"0A61", x"0A2E", x"092A", x"074C", x"0453", x"01F7", x"0133", x"0166", x"023E", x"03BF", x"04B6", x"04E5", x"0525", x"0585", x"05E5", x"0689", x"0751", x"07AE", x"080D", x"0899", x"08F5", x"0902", x"0856", x"06A3", x"040E", x"00F9", x"FDAD", x"FAD3", x"F8EE", x"F7C3", x"F7BE", x"F8E5", x"FA18", x"FB07", x"FCA1", x"FEA8", x"004C", x"01E0", x"02F6", x"0227", x"00A5", x"0068", x"012D", x"0285", x"04D5", x"06FF", x"076A", x"06BA", x"0567", x"02C6", x"FFBD", x"FDA1", x"FC52", x"FBE6", x"FCE7", x"FE71", x"FFB1", x"00FB", x"01FA", x"0212", x"0229", x"0276", x"022E", x"01C1", x"01B1", x"0150", x"00F3", x"0198", x"0270", x"0307", x"03F9", x"04F2", x"055A", x"065D", x"082E", x"09D3", x"0BB4", x"0E2C", x"0FB3", x"10B2", x"12AC", x"14A6", x"154C", x"154A", x"13E6", x"1028", x"0C7D", x"0B28", x"0B1B", x"0BE0", x"0E09", x"0FCE", x"0FCB", x"0F48", x"0E61", x"0BFE", x"0968", x"080F", x"0791", x"080A", x"09EE", x"0BC7", x"0C87", x"0CA5", x"0BF0", x"0A39", x"08A4", x"073F", x"0589", x"03EC", x"02C8", x"01B2", x"0136", x"01D0", x"029F", x"0385", x"04BF", x"05CE", x"06A4", x"081B", x"09AF", x"0AF4", x"0C73", x"0D9F", x"0D5F", x"0D04", x"0D60", x"0D7E", x"0D98", x"0DF2", x"0CD5", x"09F0", x"07DD", x"072A", x"0713", x"085B", x"0A9B", x"0B7F", x"0B37", x"0AD0", x"0971", x"0712", x"0543", x"03B5", x"0203", x"0121", x"00B1", x"FF61", x"FDD7", x"FC36", x"F9CE", x"F7C5", x"F74B", x"F769", x"F7A7", x"F89C", x"F8F7", x"F842", x"F856", x"F95B", x"FA47", x"FBE2", x"FE11", x"FF2F", x"002D", x"0247", x"0492", x"06E6", x"0A4C", x"0D02", x"0DEC", x"0F1B", x"10BA", x"115F", x"11EA", x"1271", x"109D", x"0D84", x"0C49", x"0C86", x"0D69", x"100E", x"12F3", x"139B", x"1305", x"1220", x"0F84", x"0BF5", x"0976", x"07B3", x"06B6", x"07AF", x"098C", x"0AAA", x"0B7C", x"0BD2", x"0B15", x"0A8D", x"0ADB", x"0AFF", x"0B03", x"0B17", x"0A26", x"0853", x"06C7", x"04FA", x"0292", x"0067", x"FE08", x"FB01", x"F89B", x"F759", x"F674", x"F6F4", x"F8CE", x"FA37", x"FB5D", x"FD85", x"FFCD", x"01D9", x"04C6", x"0711", x"070B", x"06B1", x"0779", x"0870", x"0A22", x"0D0B", x"0EBB", x"0E4C", x"0D39", x"0B45", x"07FD", x"04FC", x"0305", x"015E", x"00FE", x"022C", x"0382", x"04CF", x"0678", x"0744", x"0756", x"07E2", x"0853", x"081E", x"0840", x"0815", x"0682", x"051A", x"04B4", x"0449", x"0476", x"05C1", x"063A", x"05C0", x"05DA", x"0615", x"05DD", x"06E2", x"0880", x"08ED", x"09A6", x"0BD7", x"0DD3", x"0F70", x"114B", x"10D1", x"0D2E", x"0996", x"0740", x"0562", x"0548", x"06F7", x"07C2", x"075D", x"0745", x"065C", x"0412", x"0224", x"011A", x"0081", x"0177", x"03F3", x"063B", x"0804", x"0975", x"09D1", x"099F", x"09D2", x"09CB", x"0932", x"086C", x"06C6", x"03E7", x"0153", x"FF87", x"FE04", x"FD86", x"FDD3", x"FD8E", x"FD04", x"FD06", x"FCFC", x"FD04", x"FE18", x"FF0B", x"FF0E", x"FF77", x"0079", x"012A", x"026E", x"0414", x"0420", x"02EA", x"0284", x"02D1", x"0391", x"05E0", x"08A3", x"09F9", x"0A74", x"0A78", x"0909", x"06A7", x"049E", x"02B3", x"011D", x"009C", x"006A", x"FFC6", x"FF48", x"FEA3", x"FDA5", x"FD78", x"FE55", x"FF53", x"00B0", x"023C", x"025F", x"0181", x"014E", x"018B", x"024B", x"047F", x"0701", x"0848", x"094A", x"0A63", x"0ABD", x"0B28", x"0C55", x"0C8E", x"0BB3", x"0BA8", x"0BBD", x"0B7F", x"0C0E", x"0C8B", x"0AFF", x"090D", x"08C6", x"095D", x"0B29", x"0EF9", x"12A9", x"145E", x"1570", x"15D0", x"143F", x"1205", x"107F", x"0F21", x"0E82", x"0FA2", x"112D", x"120E", x"12B8", x"12D8", x"1210", x"11A3", x"11BF", x"11AD", x"11A6", x"11D4", x"1158", x"10B9", x"10DB", x"10F9", x"10A6", x"1036", x"0EC8", x"0C24", x"097E", x"0725", x"04E7", x"03AA", x"0363", x"02E2", x"02B1", x"0388", x"048C", x"05AA", x"0788", x"087C", x"078C", x"06A6", x"06BA", x"0725", x"08D4", x"0BB6", x"0D63", x"0D39", x"0C63", x"0A60", x"06C6", x"0336", x"0072", x"FE23", x"FD2B", x"FDE3", x"FEDE", x"FFB6", x"0082", x"00E7", x"00F7", x"0181", x"0211", x"027A", x"030F", x"0364", x"0330", x"0388", x"0490", x"05C9", x"079A", x"09C5", x"0ABB", x"0AC2", x"0AAA", x"09F1", x"0904", x"094C", x"09E0", x"09C6", x"0A55", x"0BBF", x"0CAF", x"0DCC", x"0F20", x"0E21", x"0ADC", x"0818", x"0648", x"052F", x"0662", x"091E", x"0AA6", x"0B4A", x"0C21", x"0B93", x"0941", x"06E4", x"04A3", x"026C", x"01E9", x"033A", x"048F", x"058E", x"063E", x"05F7", x"050E", x"045E", x"0376", x"0228", x"00F1", x"FF3C", x"FD26", x"FBB6", x"FB09", x"FAC9", x"FB95", x"FCDF", x"FD60", x"FD8F", x"FDE8", x"FDC3", x"FDBF", x"FEBD", x"FF75", x"FF81", x"002A", x"0120", x"01A7", x"02A9", x"03AC", x"02B5", x"00BE", x"FFCE", x"FF8C", x"0003", x"0246", x"04C3", x"05AA", x"0615", x"0658", x"053C", x"033A", x"018B", x"FFAB", x"FDDA", x"FCEF", x"FC3D", x"FACF", x"F921", x"F742", x"F53A", x"F3C9", x"F303", x"F25B", x"F22A", x"F23E", x"F1BB", x"F13E", x"F17D", x"F1F9", x"F320", x"F590", x"F80C", x"F9D4", x"FBEA", x"FE01", x"FF85", x"0196", x"0402", x"0524", x"0590", x"066E", x"06DD", x"0725", x"0832", x"0853", x"0615", x"0392", x"01F1", x"00DE", x"01BC", x"04F1", x"07BB", x"0936", x"0A92", x"0AD5", x"0954", x"0788", x"05DA", x"03A9", x"0222", x"021F", x"0244", x"025D", x"02CB", x"02CC", x"024C", x"0228", x"01F8", x"0151", x"00D4", x"0022", x"FEC1", x"FD7D", x"FCA1", x"FB6B", x"FA5E", x"F987", x"F802", x"F62A", x"F515", x"F447", x"F3F7", x"F4FD", x"F64D", x"F6EE", x"F7C8", x"F8E0", x"F96C", x"FAA3", x"FCA6", x"FD70", x"FCF1", x"FCF5", x"FD47", x"FDF9", x"0098", x"03D4", x"0539", x"050E", x"043C", x"01C3", x"FE69", x"FBB9", x"F95F", x"F742", x"F6BB", x"F7A7", x"F8FD", x"FA9D", x"FC60", x"FD6F", x"FE16", x"FE94", x"FE9E", x"FE84", x"FE7F", x"FE2B", x"FDD0", x"FDCA", x"FDAA", x"FD8F", x"FE5C", x"FF3B", x"FFBE", x"0071", x"00B8", x"FFC1", x"FEE3", x"FE84", x"FD81", x"FC5B", x"FC27", x"FBE0", x"FBA6", x"FCFE", x"FE76", x"FDCA", x"FBE9", x"F9DE", x"F735", x"F5AA", x"F6B5", x"F848", x"F8C2", x"F924", x"F92D", x"F7E2", x"F64E", x"F50E", x"F34D", x"F1B5", x"F19B", x"F2B2", x"F47F", x"F6F8", x"F981", x"FB70", x"FCC8", x"FD23", x"FC70", x"FB54", x"F9DA", x"F84C", x"F764", x"F6E5", x"F626", x"F5E0", x"F651", x"F67C", x"F6A1", x"F730", x"F6F5", x"F5F9", x"F5BA", x"F5C1", x"F507", x"F482", x"F460", x"F39B", x"F35A", x"F4C4", x"F5C6", x"F565", x"F4D6", x"F441", x"F3B1", x"F50D", x"F86A", x"FB4E", x"FCFA", x"FDDA", x"FD42", x"FB25", x"F8EE", x"F6CA", x"F47C", x"F2D4", x"F207", x"F191", x"F145", x"F12F", x"F115", x"F14C", x"F1A5", x"F1A7", x"F1A9", x"F1E8", x"F20F", x"F287", x"F3B4", x"F490", x"F4F4", x"F5E7", x"F720", x"F81C", x"F9C6", x"FBAD", x"FC9D", x"FD16", x"FDEF", x"FDD5", x"FCDA", x"FC34", x"FB72", x"FA8C", x"FB4E", x"FD82", x"FED4", x"FF3A", x"FF0D", x"FDB2", x"FC53", x"FD03", x"FEF9", x"00A7", x"0252", x"0386", x"0349", x"025C", x"0189", x"0044", x"FEF2", x"FE75", x"FE90", x"FF4A", x"00D2", x"02D9", x"04CB", x"06C3", x"07F6", x"07F6", x"0774", x"0694", x"0575", x"04F1", x"04F4", x"0469", x"038F", x"02C0", x"014A", x"FF67", x"FE1D", x"FC61", x"F9D9", x"F7C4", x"F63A", x"F471", x"F38D", x"F3F3", x"F434", x"F4E2", x"F720", x"F968", x"FA4E", x"FAA7", x"FA33", x"F89E", x"F815", x"F9BE", x"FBAF", x"FCD6", x"FD5B", x"FC34", x"F95A", x"F66F", x"F3FA", x"F174", x"EF89", x"EEB7", x"EEA6", x"EF56", x"F0D7", x"F28F", x"F41D", x"F56E", x"F621", x"F678", x"F701", x"F7A2", x"F8FF", x"FB5B", x"FDC7", x"FF6C", x"00BA", x"0144", x"00F4", x"0135", x"0245", x"02C8", x"02FB", x"038E", x"035F", x"0282", x"0258", x"0241", x"0160", x"0159", x"02A2", x"0353", x"02E6", x"01F4", x"FF62", x"FBEA", x"FA38", x"FAC4", x"FBEF", x"FD99", x"FF52", x"FFF0", x"FF75", x"FEF5", x"FDD9", x"FBDB", x"F99B", x"F793", x"F5D8", x"F4CA", x"F46E", x"F496", x"F51B", x"F56D", x"F50F", x"F423", x"F287", x"F071", x"EF1D", x"EED8", x"EEA4", x"EE85", x"EECD", x"EEB5", x"EEA0", x"EFD6", x"F196", x"F294", x"F399", x"F4EB", x"F562", x"F5A9", x"F69B", x"F6F0", x"F664", x"F6F6", x"F880", x"F947", x"F995", x"F984", x"F833", x"F6F9", x"F823", x"FB22", x"FE11", x"00AA", x"020C", x"00FD", x"FE4D", x"FB13", x"F73E", x"F2F5", x"EF75", x"ECF2", x"EB3B", x"EA59", x"EA0D", x"E9C3", x"E96A", x"E8B5", x"E7CC", x"E6C9", x"E5F9", x"E5AD", x"E678", x"E801", x"E94E", x"EA4A", x"EAC0", x"EA7B", x"EA4D", x"EB53", x"ECFC", x"EEC0", x"F119", x"F35F", x"F487", x"F547", x"F608", x"F5EF", x"F5C5", x"F711", x"F8EA", x"FA20", x"FAFC", x"FB2C", x"FA0E", x"F98E", x"FB25", x"FDBF", x"004C", x"02C9", x"0410", x"0375", x"020C", x"0056", x"FDCD", x"FB0A", x"F8E2", x"F73F", x"F657", x"F6A1", x"F7AF", x"F8F0", x"FA45", x"FB1B", x"FB02", x"FA69", x"F96B", x"F870", x"F81A", x"F829", x"F7FC", x"F7A1", x"F710", x"F5FC", x"F56F", x"F5FD", x"F6B4", x"F742", x"F813", x"F82E", x"F72D", x"F688", x"F62E", x"F549", x"F540", x"F707", x"F8C9", x"F9E5", x"FAF0", x"FACA", x"F959", x"F999", x"FC15", x"FEE3", x"0149", x"030E", x"0243", x"FF55", x"FCA7", x"FA2C", x"F766", x"F594", x"F52A", x"F563", x"F6E0", x"F9F2", x"FCF1", x"FF23", x"00B8", x"013B", x"0088", x"FFAF", x"FEE8", x"FE32", x"FE2D", x"FEC6", x"FF65", x"000A", x"0062", x"003A", x"0068", x"0128", x"01D0", x"0284", x"033C", x"02D7", x"0181", x"0066", x"FEE6", x"FCE5", x"FC65", x"FD7E", x"FE86", x"FF5A", x"FFE6", x"FE44", x"FB7B", x"FA5D", x"FAD8", x"FB8F", x"FCEA", x"FE21", x"FD9C", x"FC64", x"FBE4", x"FB2F", x"F9F7", x"F979", x"F976", x"F998", x"FAA8", x"FC7F", x"FDE4", x"FEEA", x"FF91", x"FF5A", x"FE7F", x"FD6A", x"FC21", x"FB2D", x"FADF", x"FAC5", x"FAB6", x"FABF", x"FA45", x"F9B0", x"FA09", x"FAB3", x"FB0F", x"FBE8", x"FCBD", x"FC7D", x"FC14", x"FC1C", x"FAE5", x"F931", x"F949", x"FA5C", x"FB21", x"FC71", x"FD2F", x"FBAE", x"FA41", x"FB64", x"FDBE", x"004D", x"0369", x"0520", x"043D", x"02EA", x"020A", x"0067", x"FE9D", x"FDC6", x"FCE3", x"FC20", x"FC9F", x"FD7A", x"FD9D", x"FD8D", x"FD19", x"FBC0", x"FA7C", x"F9EA", x"F9BB", x"FA47", x"FBCB", x"FD34", x"FE54", x"FF2D", x"FF49", x"FF19", x"FFB9", x"00F2", x"027B", x"04D3", x"06F3", x"07B9", x"081A", x"0843", x"0778", x"0739", x"08D6", x"0AE2", x"0C2D", x"0D32", x"0C55", x"0927", x"06A3", x"0685", x"079C", x"09E5", x"0D34", x"0F47", x"0FA2", x"1002", x"102F", x"0F5A", x"0E97", x"0E3F", x"0D95", x"0D5D", x"0E5E", x"0F85", x"1093", x"11D4", x"126B", x"1223", x"11BC", x"1129", x"1076", x"1047", x"107E", x"1056", x"1016", x"0F4B", x"0D76", x"0B88", x"09F3", x"0827", x"069F", x"05CB", x"045B", x"029E", x"01C4", x"00F6", x"FF98", x"FFC1", x"0170", x"02EF", x"04AB", x"0663", x"059A", x"031C", x"024F", x"0327", x"049E", x"0746", x"0986", x"089D", x"0611", x"03D0", x"010E", x"FE11", x"FC76", x"FB51", x"FA1D", x"FA95", x"FC7C", x"FE3F", x"0041", x"02A9", x"0451", x"05C4", x"07E1", x"09B6", x"0AF3", x"0C28", x"0CE0", x"0CB2", x"0C71", x"0BD8", x"0ABC", x"0A16", x"0A31", x"0A6C", x"0B68", x"0CA6", x"0CDE", x"0C7A", x"0C23", x"0AAB", x"08BC", x"0848", x"08CD", x"0945", x"0A57", x"0AA1", x"0807", x"0478", x"028C", x"01DE", x"027C", x"0506", x"0741", x"0774", x"0730", x"06D9", x"054D", x"033B", x"017B", x"FF57", x"FD3D", x"FC91", x"FCD9", x"FDA1", x"FF36", x"011B", x"024A", x"02D4", x"0285", x"0131", x"FFB3", x"FE76", x"FD78", x"FCE5", x"FC93", x"FBD4", x"FB6A", x"FBF0", x"FCD5", x"FE3C", x"00A8", x"02A0", x"03A7", x"04F7", x"05C0", x"04E1", x"03FD", x"0444", x"04AD", x"05A7", x"0806", x"093C", x"086C", x"0855", x"09FF", x"0C66", x"100B", x"1426", x"1573", x"139A", x"10C6", x"0D0A", x"0882", x"04F6", x"0282", x"000C", x"FE5F", x"FDFA", x"FD96", x"FD14", x"FCCE", x"FBF2", x"FA32", x"F87C", x"F6D5", x"F55A", x"F4C9", x"F532", x"F5DA", x"F6CD", x"F7A3", x"F7E2", x"F838", x"F95C", x"FB38", x"FE18", x"01D8", x"04B1", x"0607", x"0644", x"04E5", x"021C", x"0020", x"FFA6", x"FFE4", x"0144", x"0354", x"03DA", x"02CE", x"02AA", x"03D1", x"060B", x"0A24", x"0EF0", x"1202", x"1356", x"140D", x"1379", x"11D1", x"106E", x"0F46", x"0DEF", x"0D55", x"0D9D", x"0DE7", x"0E38", x"0EB7", x"0EC0", x"0E1E", x"0D15", x"0B7B", x"097C", x"07C0", x"0680", x"05DF", x"05CB", x"05A5", x"0524", x"04B7", x"0417", x"036C", x"0323", x"02A6", x"010E", x"FF4F", x"FDE7", x"FC1E", x"FAA4", x"FAE8", x"FBEE", x"FD54", x"FFE8", x"0251", x"0251", x"0164", x"0168", x"020D", x"03BF", x"0720", x"0973", x"08B3", x"065F", x"036B", x"FF88", x"FC36", x"FAC5", x"F9E3", x"F9BA", x"FB56", x"FDC0", x"FFBE", x"01BA", x"0364", x"03F6", x"0451", x"0531", x"05E0", x"06B8", x"0833", x"09E2", x"0B92", x"0D62", x"0E94", x"0ECC", x"0EAE", x"0E64", x"0E1A", x"0E6C", x"0E92", x"0DA0", x"0C14", x"09DB", x"065D", x"02EF", x"0108", x"FFFA", x"FFD8", x"0102", x"013D", x"FF00", x"FC33", x"FA78", x"F98D", x"FA92", x"FDAC", x"002A", x"0124", x"0220", x"0315", x"032F", x"0362", x"03C3", x"02EB", x"018A", x"009C", x"FFA8", x"FE8C", x"FE57", x"FEA8", x"FEE0", x"FF2B", x"FF0A", x"FE10", x"FCC5", x"FBDF", x"FB79", x"FBBF", x"FC43", x"FC64", x"FC5E", x"FC88", x"FCE5", x"FE19", x"0023", x"01B0", x"02AD", x"0399", x"0381", x"0225", x"013E", x"011F", x"0104", x"020E", x"03E4", x"03B4", x"015A", x"FF44", x"FDEA", x"FD96", x"0002", x"03CF", x"05CD", x"063F", x"064E", x"0525", x"034D", x"0288", x"020A", x"0102", x"00EC", x"01C2", x"0241", x"02CC", x"03B3", x"03A7", x"02EC", x"028B", x"022C", x"01BE", x"023F", x"0332", x"03D9", x"0474", x"04B2", x"03F3", x"02FD", x"028B", x"028E", x"03DB", x"0666", x"08C3", x"0A81", x"0B9B", x"0AF1", x"08B6", x"0707", x"05FB", x"0543", x"0601", x"0733", x"064E", x"042B", x"02F8", x"0296", x"03A0", x"0799", x"0C35", x"0F04", x"10E4", x"127F", x"1271", x"11E5", x"11F3", x"1160", x"1019", x"0FD2", x"102C", x"1037", x"10E6", x"1210", x"129B", x"1324", x"142A", x"14B1", x"14C6", x"14D6", x"145C", x"1337", x"1226", x"10BB", x"0EF0", x"0D85", x"0C7E", x"0BCD", x"0C36", x"0CCA", x"0C7D", x"0BF1", x"0AF5", x"087F", x"05FA", x"04D1", x"03FD", x"03FD", x"05EF", x"0747", x"05ED", x"03FB", x"02B0", x"018D", x"02D0", x"06CE", x"0971", x"0939", x"07CD", x"04DF", x"0055", x"FD25", x"FB59", x"F916", x"F7B0", x"F84C", x"F97F", x"FB65", x"FEFD", x"0255", x"0498", x"0714", x"0947", x"0A61", x"0BA3", x"0D0E", x"0D6B", x"0DB6", x"0E74", x"0E72", x"0E47", x"0ED1", x"0F0C", x"0F3D", x"1081", x"115E", x"1132", x"1116", x"1015", x"0CEA", x"09D9", x"07BE", x"0580", x"04CA", x"0632", x"0630", x"03D8", x"01DA", x"0067", x"FFA6", x"0267", x"0765", x"0A53", x"0B51", x"0B8C", x"09C9", x"06E7", x"053A", x"033A", x"FFD7", x"FD27", x"FB5F", x"F989", x"F944", x"FA98", x"FB90", x"FC61", x"FD7F", x"FD73", x"FC8D", x"FC23", x"FB57", x"F9E4", x"F934", x"F897", x"F798", x"F79E", x"F8AE", x"F979", x"FB1C", x"FD60", x"FE6F", x"FF11", x"0035", x"FFD3", x"FE41", x"FD92", x"FD21", x"FCC6", x"FF37", x"031D", x"04C8", x"0503", x"0513", x"03B8", x"031D", x"05C4", x"089D", x"0918", x"08A0", x"06D3", x"02A2", x"FF06", x"FCDE", x"F9F1", x"F6E9", x"F554", x"F3B7", x"F231", x"F275", x"F2CD", x"F19B", x"F060", x"EED6", x"EC2B", x"EA79", x"EA74", x"EA2C", x"E9FF", x"EAC1", x"EAEA", x"EAF6", x"ECA0", x"EED1", x"F0CF", x"F3DF", x"F6D7", x"F836", x"F980", x"FA7D", x"F945", x"F77F", x"F6B5", x"F59F", x"F576", x"F84D", x"FB2F", x"FBA9", x"FBB4", x"FB6F", x"FA65", x"FC1D", x"019F", x"06C4", x"0A4E", x"0D2D", x"0DA3", x"0BD6", x"0AFC", x"0A90", x"08AB", x"06D2", x"057C", x"0328", x"0147", x"0118", x"00A4", x"FFA8", x"FF64", x"FEC1", x"FD99", x"FDDE", x"FEE6", x"FF3F", x"FFB0", x"0018", x"FF12", x"FE1E", x"FE12", x"FD99", x"FD45", x"FDC4", x"FD4C", x"FBC0", x"FAFA", x"F999", x"F6EF", x"F523", x"F41A", x"F273", x"F2C1", x"F5B7", x"F76E", x"F749", x"F704", x"F555", x"F31D", x"F496", x"F887", x"FAFB", x"FC26", x"FC3D", x"F964", x"F5E5", x"F4C9", x"F439", x"F351", x"F3A7", x"F40F", x"F374", x"F3F5", x"F58B", x"F62A", x"F6FC", x"F874", x"F91B", x"FA03", x"FCC7", x"FF6D", x"0166", x"03C6", x"053D", x"0526", x"05F3", x"0749", x"07A0", x"0847", x"0905", x"07B0", x"05BB", x"04D6", x"02CE", x"FFD5", x"FE12", x"FBC1", x"F86E", x"F765", x"F7EB", x"F665", x"F410", x"F1FC", x"EE89", x"EC45", x"EEAF", x"F2E9", x"F613", x"F926", x"FABF", x"F936", x"F792", x"F6EC", x"F510", x"F2C3", x"F150", x"EF2B", x"ECF8", x"ECFD", x"EDE1", x"EEA1", x"F06A", x"F1F1", x"F1A7", x"F1B7", x"F26D", x"F1E0", x"F116", x"F0B6", x"EEE0", x"EC9E", x"EC64", x"ECBD", x"ED01", x"EEE7", x"F0C0", x"F12E", x"F264", x"F47B", x"F4F4", x"F53F", x"F628", x"F589", x"F4AE", x"F65F", x"F82A", x"F7FF", x"F7B6", x"F6A2", x"F3E4", x"F36B", x"F69E", x"F9F9", x"FCA0", x"FEF8", x"FEAB", x"FC07", x"FA69", x"F952", x"F769", x"F669", x"F5BE", x"F3E3", x"F29F", x"F2F1", x"F2CC", x"F28B", x"F305", x"F20F", x"F008", x"EF6A", x"EF68", x"EEC2", x"EF10", x"EFA5", x"EEE7", x"EF08", x"F128", x"F369", x"F634", x"FA58", x"FD66", x"FEFB", x"00E6", x"01AB", x"003C", x"FEBF", x"FD14", x"F9E9", x"F80D", x"F88B", x"F85B", x"F742", x"F679", x"F459", x"F1BE", x"F2DB", x"F720", x"FB84", x"001E", x"040B", x"04A5", x"03CD", x"0408", x"03D8", x"031C", x"0349", x"0332", x"0208", x"0243", x"03BD", x"04DF", x"06A3", x"08E5", x"098F", x"0999", x"0A7A", x"0A69", x"0925", x"07E1", x"059D", x"01FD", x"FFAC", x"FECE", x"FE15", x"FE75", x"FFB2", x"FF9A", x"FF07", x"FF3E", x"FE6D", x"FCC7", x"FBEE", x"FA7F", x"F82F", x"F7F5", x"F992", x"FA2A", x"FA78", x"FAA6", x"F89B", x"F67F", x"F7BB", x"FA54", x"FBCD", x"FCEF", x"FC23", x"F7FA", x"F374", x"F07D", x"ED72", x"EAF9", x"EA50", x"E9CB", x"E934", x"EA57", x"EC1D", x"ED91", x"EFFC", x"F2C9", x"F49B", x"F6F1", x"FA1C", x"FC5F", x"FE35", x"0055", x"010A", x"010E", x"0268", x"0419", x"052A", x"06E4", x"07F0", x"06C8", x"057D", x"04B1", x"0281", x"0031", x"FECB", x"FC47", x"F971", x"F951", x"FA00", x"F965", x"F904", x"F84B", x"F5BE", x"F4FB", x"F838", x"FC31", x"FF7D", x"02C0", x"0382", x"0150", x"FF85", x"FE59", x"FC25", x"FA58", x"F94C", x"F747", x"F582", x"F57A", x"F5A2", x"F62A", x"F7E6", x"F8B3", x"F7F1", x"F77B", x"F6D3", x"F4F1", x"F3BE", x"F2F7", x"F0C5", x"EF4A", x"F008", x"F0D4", x"F1CD", x"F42C", x"F5AE", x"F5E4", x"F798", x"FA07", x"FB12", x"FCAB", x"FEC5", x"FF54", x"0090", x"0475", x"07B9", x"0921", x"0A25", x"091A", x"05E5", x"0508", x"0700", x"089F", x"0A03", x"0B1E", x"0939", x"05A4", x"0346", x"00F5", x"FDFB", x"FBFC", x"FA14", x"F71B", x"F53B", x"F492", x"F3A0", x"F371", x"F3FD", x"F317", x"F1AD", x"F192", x"F13A", x"F08E", x"F13B", x"F19E", x"F0CA", x"F1A6", x"F42F", x"F623", x"F861", x"FB02", x"FB58", x"FA89", x"FACE", x"FA60", x"F8B5", x"F7DE", x"F6A3", x"F423", x"F37D", x"F506", x"F5E3", x"F6B4", x"F7D9", x"F6FA", x"F5CF", x"F842", x"FCFF", x"0212", x"0830", x"0D4B", x"0EE4", x"0F6B", x"105B", x"0FDD", x"0EA7", x"0E0D", x"0C39", x"0989", x"0856", x"07C7", x"06FA", x"0784", x"0840", x"0760", x"06C4", x"06F1", x"05D7", x"0460", x"036E", x"00D8", x"FD5D", x"FC10", x"FBD5", x"FB86", x"FCC9", x"FE4E", x"FDE9", x"FDDC", x"FF15", x"FF1B", x"FEC2", x"FF16", x"FDD8", x"FB7D", x"FBA7", x"FCF4", x"FD53", x"FE29", x"FE47", x"FB69", x"F91E", x"FA73", x"FCB1", x"FF1B", x"0247", x"032F", x"00DA", x"FF18", x"FE69", x"FCD7", x"FC0D", x"FC43", x"FB49", x"FA30", x"FABA", x"FB3D", x"FBE7", x"FE40", x"00C2", x"0282", x"0559", x"086B", x"0A43", x"0C94", x"0EFA", x"0F66", x"0F85", x"10DB", x"1159", x"115A", x"124F", x"11BF", x"0F18", x"0D4F", x"0BD0", x"08CE", x"0677", x"0488", x"0066", x"FCAA", x"FBB1", x"FAF1", x"F9B7", x"F9C2", x"F899", x"F5AE", x"F5D7", x"F9CC", x"FE45", x"0367", x"0889", x"09BB", x"082D", x"0712", x"056B", x"0271", x"0063", x"FE5B", x"FB31", x"F94C", x"F91F", x"F93A", x"FACB", x"FDD6", x"FF93", x"006C", x"0187", x"0125", x"FFEB", x"FFEE", x"FF36", x"FCE7", x"FC21", x"FCE7", x"FD5D", x"FF95", x"033A", x"04A7", x"0552", x"07C4", x"09C3", x"0A9F", x"0CA2", x"0D2E", x"0A8D", x"08DF", x"0905", x"0812", x"0739", x"06F6", x"03F7", x"FFB2", x"FEDF", x"0041", x"01E8", x"051F", x"07DA", x"072E", x"05B9", x"054B", x"03ED", x"026D", x"0234", x"015D", x"000D", x"0041", x"010F", x"0186", x"0344", x"04D0", x"0483", x"041C", x"03E2", x"0267", x"018A", x"0208", x"012D", x"FFE6", x"00B3", x"020B", x"0341", x"062F", x"0894", x"0804", x"074A", x"0785", x"069C", x"0612", x"06E8", x"05FB", x"03B1", x"0388", x"0459", x"049B", x"0602", x"0704", x"04F5", x"0309", x"0402", x"0633", x"09D4", x"0F70", x"1381", x"149A", x"1558", x"15A1", x"14B3", x"1468", x"14DA", x"1427", x"1399", x"1439", x"14AC", x"15BB", x"1848", x"1A0C", x"1A67", x"1ACE", x"1A14", x"17FD", x"16DD", x"160A", x"1392", x"117B", x"10B8", x"0F8F", x"0F3C", x"1124", x"1222", x"119F", x"11FF", x"1220", x"1097", x"0FC3", x"0EF4", x"0B85", x"07E5", x"069A", x"056E", x"046B", x"04D6", x"0383", x"FF66", x"FCBA", x"FCD5", x"FDD3", x"00C8", x"04DF", x"061B", x"04F1", x"043E", x"0349", x"01CF", x"01B6", x"01E9", x"00C6", x"0020", x"0047", x"0029", x"00F4", x"035A", x"058E", x"07E2", x"0B11", x"0D96", x"0F9F", x"12AB", x"1552", x"16AA", x"1883", x"1A57", x"1AF6", x"1C3E", x"1E10", x"1DBE", x"1C26", x"1AF0", x"1882", x"1564", x"1403", x"127B", x"0F38", x"0D5B", x"0D3B", x"0C9E", x"0C99", x"0D5D", x"0B8B", x"0807", x"06DA", x"0783", x"08B1", x"0B9C", x"0E45", x"0DA6", x"0BA3", x"09FA", x"075C", x"046B", x"02AB", x"00B0", x"FE68", x"FD8F", x"FD7A", x"FD86", x"FEC6", x"007C", x"013B", x"01EC", x"024D", x"0141", x"0057", x"0027", x"FECD", x"FCDB", x"FBFD", x"FADD", x"F9EC", x"FB72", x"FD69", x"FD89", x"FDFA", x"FF04", x"FEF1", x"FFD6", x"02AC", x"03CD", x"0314", x"03F8", x"0567", x"063D", x"0895", x"0AEA", x"09AA", x"07A3", x"0803", x"0926", x"0B49", x"0F59", x"122B", x"11A3", x"107F", x"0F17", x"0C1F", x"094F", x"072A", x"0402", x"00A3", x"FE64", x"FC2E", x"FA2C", x"F9AB", x"F951", x"F882", x"F855", x"F7F1", x"F6B9", x"F676", x"F6B9", x"F5FD", x"F586", x"F5FC", x"F5D9", x"F64F", x"F89C", x"FA19", x"FA25", x"FACE", x"FB40", x"FA9A", x"FB5A", x"FCE8", x"FC46", x"FB1D", x"FB97", x"FBD7", x"FBFC", x"FD81", x"FDAA", x"FAF3", x"F922", x"F9F4", x"FC39", x"0102", x"07D4", x"0CB7", x"0EED", x"1029", x"0FEB", x"0E2C", x"0D1B", x"0C7D", x"0B62", x"0B07", x"0B80", x"0BD1", x"0CD8", x"0EBC", x"0FDF", x"1042", x"1040", x"0E9E", x"0C2F", x"0A94", x"08E7", x"06B1", x"0563", x"0448", x"029D", x"029A", x"044B", x"055B", x"065A", x"0817", x"0853", x"079E", x"0845", x"084F", x"0634", x"04CB", x"0489", x"037A", x"0332", x"0410", x"025C", x"FE9C", x"FCB2", x"FCAF", x"FDC6", x"0183", x"05EA", x"0739", x"0698", x"059C", x"0333", x"001E", x"FE28", x"FC09", x"F945", x"F7B2", x"F6F3", x"F635", x"F6CD", x"F89C", x"FA84", x"FD3B", x"0114", x"047C", x"07E1", x"0BBA", x"0E93", x"1068", x"1294", x"1427", x"1512", x"1709", x"18DB", x"18B9", x"17AB", x"15D8", x"11CE", x"0DA9", x"0B21", x"07E2", x"03D1", x"0190", x"0021", x"FE4D", x"FE07", x"FE1F", x"FB49", x"F785", x"F618", x"F616", x"F7BF", x"FC4D", x"00C3", x"028D", x"0377", x"03FE", x"02B7", x"0101", x"FFD1", x"FDEF", x"FBFF", x"FB8A", x"FB8E", x"FBD2", x"FD1D", x"FE84", x"FF31", x"0006", x"005A", x"FF4A", x"FE25", x"FCB6", x"FA33", x"F7B1", x"F620", x"F47C", x"F411", x"F631", x"F891", x"FA72", x"FCF8", x"FE97", x"FEA1", x"FFB4", x"0179", x"010C", x"FFFF", x"0039", x"0004", x"0011", x"026B", x"03B5", x"0186", x"FF1D", x"FE18", x"FD58", x"FEAD", x"0242", x"0407", x"031D", x"01FA", x"000A", x"FD36", x"FBA1", x"FAE8", x"F95D", x"F80E", x"F750", x"F5D8", x"F491", x"F490", x"F48B", x"F4E7", x"F67E", x"F819", x"F970", x"FBAF", x"FDCF", x"FEEB", x"0047", x"0192", x"01F4", x"030F", x"0537", x"066F", x"0714", x"07EE", x"0712", x"0542", x"04CA", x"0443", x"0221", x"00D6", x"009C", x"FFCD", x"0026", x"0204", x"01A8", x"FEB6", x"FC9E", x"FBB7", x"FBE5", x"FF46", x"046A", x"0798", x"093A", x"0A70", x"0A5A", x"09A9", x"0A2C", x"0B18", x"0BCB", x"0D58", x"0F02", x"0FDD", x"10B8", x"1167", x"1103", x"1046", x"0F46", x"0D22", x"0AC6", x"08D7", x"0693", x"043B", x"02C2", x"0133", x"FFD2", x"0028", x"0176", x"02AE", x"04A8", x"0687", x"06A8", x"06D4", x"080F", x"0838", x"0757", x"071D", x"0615", x"03C4", x"0298", x"01A5", x"FDFE", x"F984", x"F6B7", x"F4F8", x"F52A", x"F884", x"FC12", x"FCEB", x"FC60", x"FABF", x"F754", x"F3B3", x"F120", x"EE97", x"EC79", x"EBCD", x"EBB1", x"EBD5", x"ED30", x"EF4F", x"F1C1", x"F554", x"F98D", x"FD53", x"010C", x"046B", x"066B", x"07A1", x"08B9", x"090A", x"091D", x"09D4", x"09FD", x"092E", x"082A", x"0607", x"0262", x"FF66", x"FD52", x"FAAB", x"F86D", x"F7A8", x"F6A0", x"F5EA", x"F6E3", x"F74A", x"F4CD", x"F1D4", x"EFDF", x"EE9E", x"EFCA", x"F405", x"F802", x"FA1B", x"FB9C", x"FC09", x"FAB4", x"F905", x"F778", x"F505", x"F297", x"F0E4", x"EF30", x"EDAA", x"ED0F", x"ECAF", x"EC6B", x"ECB7", x"ECBE", x"EBF8", x"EAF8", x"E989", x"E74A", x"E581", x"E496", x"E441", x"E55C", x"E815", x"EB3A", x"EEBC", x"F2A8", x"F567", x"F713", x"F91F", x"FAAE", x"FAF5", x"FBAA", x"FCC9", x"FD45", x"FEB9", x"01A6", x"02DE", x"018B", x"0003", x"FE7F", x"FD4B", x"FEB6", x"01E0", x"0356", x"02DB", x"018E", x"FE9D", x"FAAA", x"F7A6", x"F4F3", x"F1E1", x"EF50", x"ED09", x"EA45", x"E813", x"E718", x"E6C8", x"E7B4", x"EA1A", x"ECAC", x"EEF2", x"F12C", x"F224", x"F196", x"F073", x"EEDC", x"ECA8", x"EB1F", x"EA3A", x"E976", x"E95C", x"E99D", x"E902", x"E83A", x"E817", x"E786", x"E6BD", x"E70D", x"E76E", x"E799", x"E954", x"EBE7", x"EC9B", x"EC2C", x"EC46", x"EC9E", x"EE6F", x"F373", x"F981", x"FDD9", x"00ED", x"0303", x"035B", x"0325", x"03BB", x"0459", x"04DE", x"05F5", x"06D0", x"06AB", x"0621", x"0527", x"038C", x"0215", x"00C5", x"FF17", x"FD50", x"FBA7", x"F9B2", x"F7F3", x"F706", x"F6AE", x"F6F5", x"F7FF", x"F954", x"FAB3", x"FC76", x"FDAB", x"FDE5", x"FDF6", x"FDE0", x"FCF4", x"FC22", x"FB9E", x"FA2B", x"F85E", x"F7A5", x"F669", x"F374", x"F04B", x"EDFE", x"EC64", x"ED14", x"F093", x"F3E7", x"F547", x"F588", x"F4AD", x"F26B", x"F044", x"EF10", x"EE0B", x"ED7D", x"EDFA", x"EEB2", x"EF2B", x"F004", x"F13F", x"F2D5", x"F55B", x"F86B", x"FB58", x"FE05", x"004A", x"01C1", x"02E8", x"045F", x"05D4", x"072D", x"084F", x"08BA", x"084B", x"0772", x"05DF", x"039E", x"0180", x"FF46", x"FCD7", x"FAFE", x"F9FB", x"F906", x"F8F0", x"F9FE", x"FA06", x"F7D6", x"F4F4", x"F21B", x"EFEF", x"F08F", x"F434", x"F7F9", x"FABB", x"FD1E", x"FE3A", x"FD92", x"FC65", x"FAEB", x"F877", x"F5F2", x"F419", x"F24E", x"F0A4", x"EFD1", x"EF66", x"EF52", x"EFEE", x"F07B", x"F092", x"F080", x"F007", x"EED1", x"EDDD", x"EDCB", x"EE51", x"EFB9", x"F20D", x"F457", x"F681", x"F8D0", x"FA98", x"FBA2", x"FC59", x"FC27", x"FAF6", x"F9E6", x"F90B", x"F830", x"F883", x"F9BD", x"F981", x"F7A0", x"F54B", x"F2B9", x"F0E4", x"F206", x"F4F6", x"F713", x"F850", x"F8FB", x"F837", x"F6D6", x"F665", x"F630", x"F5D5", x"F5EC", x"F61B", x"F56D", x"F4DB", x"F4C0", x"F4EA", x"F622", x"F87E", x"FB12", x"FD9E", x"0027", x"017D", x"0150", x"00B1", x"FFA9", x"FE4E", x"FD80", x"FD44", x"FD0A", x"FD59", x"FE31", x"FED1", x"FF2C", x"FF53", x"FEA4", x"FDB9", x"FD70", x"FD2F", x"FD54", x"FEB5", x"0012", x"FFAC", x"FE1E", x"FBF3", x"F92D", x"F803", x"F9FF", x"FD30", x"0002", x"02A6", x"0481", x"04F3", x"0582", x"06E6", x"0836", x"09B6", x"0BCA", x"0D8A", x"0E95", x"0F76", x"1006", x"1010", x"105C", x"108D", x"1024", x"0F72", x"0E56", x"0C74", x"0A52", x"08DF", x"07F2", x"079E", x"0810", x"0894", x"08FF", x"09BC", x"0A9C", x"0B6C", x"0C5E", x"0D10", x"0D04", x"0CDC", x"0C70", x"0B11", x"09A0", x"08B4", x"0700", x"040D", x"00FD", x"FE01", x"FB95", x"FBF7", x"FF28", x"029A", x"04F5", x"066E", x"0626", x"043C", x"025A", x"00DA", x"FF04", x"FD99", x"FD2A", x"FD08", x"FD0A", x"FDC9", x"FF1D", x"0114", x"0417", x"07B2", x"0B3F", x"0E87", x"112D", x"12E2", x"1430", x"155B", x"1631", x"16F0", x"175B", x"1714", x"1644", x"1557", x"1413", x"12A9", x"1162", x"0FA4", x"0D53", x"0B42", x"0944", x"0772", x"0707", x"07F0", x"0807", x"069D", x"040C", x"000F", x"FBE2", x"FA6C", x"FB88", x"FD3F", x"FF66", x"01B4", x"02DA", x"02FE", x"0346", x"0318", x"0208", x"012A", x"009C", x"FFC8", x"FF1A", x"FED6", x"FEBA", x"FEFD", x"FFA1", x"FFC9", x"FF85", x"FF00", x"FDE6", x"FC8D", x"FBC2", x"FB3E", x"FB0F", x"FBF0", x"FD60", x"FE92", x"FFEB", x"014B", x"0205", x"0298", x"0366", x"036B", x"02FA", x"0304", x"0336", x"03F2", x"0692", x"0A12", x"0C60", x"0D77", x"0D59", x"0BA5", x"0A50", x"0B5A", x"0D87", x"0F67", x"10F3", x"113D", x"0F71", x"0CE6", x"0A93", x"080C", x"05C8", x"0423", x"0248", x"FFED", x"FD97", x"FB77", x"FA12", x"FA2A", x"FB34", x"FCC0", x"FEF4", x"012F", x"02B8", x"03D2", x"0442", x"035A", x"01DB", x"0085", x"FEE4", x"FD6D", x"FCCD", x"FC84", x"FC4A", x"FCAB", x"FCD4", x"FC26", x"FB77", x"FAF1", x"FA45", x"FA96", x"FC72", x"FE43", x"FF65", x"0001", x"FF54", x"FDBB", x"FDBE", x"0004", x"037B", x"07E1", x"0C8F", x"1008", x"1246", x"147F", x"1689", x"1855", x"1A4C", x"1C09", x"1CC3", x"1C9F", x"1BB4", x"1A06", x"1851", x"16D5", x"1524", x"136D", x"11A9", x"0F7C", x"0D20", x"0B49", x"09D4", x"08F2", x"0910", x"09C1", x"0A43", x"0ADD", x"0B50", x"0B50", x"0B5F", x"0BB2", x"0BAF", x"0B88", x"0BAF", x"0B75", x"0AB0", x"0A66", x"0A35", x"0937", x"07A0", x"057A", x"0224", x"FEDD", x"FDA9", x"FE63", x"FFFE", x"01FB", x"0346", x"029E", x"0095", x"FE46", x"FBE8", x"F9A8", x"F852", x"F7F7", x"F81A", x"F8C6", x"FA07", x"FBE9", x"FE78", x"01D2", x"05A2", x"0976", x"0CDE", x"0FC1", x"126E", x"14FC", x"174E", x"195C", x"1B04", x"1BAE", x"1B7A", x"1ADF", x"19CC", x"1880", x"177B", x"16AB", x"153B", x"1356", x"10FF", x"0DC1", x"0A3B", x"07E4", x"0651", x"04A1", x"028B", x"FFA3", x"FB60", x"F79F", x"F694", x"F830", x"FB98", x"0081", x"0593", x"093C", x"0BC5", x"0D84", x"0DE3", x"0CE8", x"0B87", x"09AE", x"0737", x"0473", x"01F0", x"FFCD", x"FE8A", x"FE21", x"FE23", x"FDF8", x"FD46", x"FC2A", x"FB37", x"FA87", x"F9FA", x"F9E4", x"FA7A", x"FB3C", x"FC95", x"FEC3", x"0117", x"033A", x"05B7", x"07F6", x"0927", x"09DC", x"0A34", x"09D2", x"09AB", x"0ACF", x"0BFE", x"0C2E", x"0B64", x"08FE", x"04FF", x"01A9", x"0068", x"008C", x"01C2", x"03C7", x"051A", x"050D", x"0470", x"0381", x"0223", x"012F", x"0114", x"0130", x"014B", x"0161", x"015E", x"01B3", x"02E6", x"04A0", x"06D3", x"0937", x"0B4A", x"0D00", x"0E9B", x"0F82", x"0F52", x"0EC4", x"0DE9", x"0C90", x"0B60", x"0AA4", x"09C1", x"08E3", x"08CC", x"087D", x"078A", x"0676", x"052A", x"03A5", x"0320", x"0409", x"0510", x"05AA", x"05A3", x"0450", x"021E", x"0103", x"018E", x"0337", x"05F0", x"0918", x"0B6F", x"0CCF", x"0E05", x"0F13", x"100E", x"1193", x"1373", x"14F8", x"15BF", x"15BE", x"14DD", x"13A3", x"1278", x"1191", x"10B8", x"0FB1", x"0E2D", x"0C70", x"0AC5", x"0934", x"084D", x"0853", x"08EC", x"09B2", x"0AC5", x"0BB8", x"0C4E", x"0D49", x"0ED8", x"1062", x"11C5", x"1317", x"1386", x"132B", x"12E0", x"127F", x"10FA", x"0E72", x"0AAE", x"053D", x"FF7A", x"FB79", x"F961", x"F8B1", x"F957", x"FA1F", x"F98A", x"F838", x"F6F2", x"F55F", x"F3EC", x"F381", x"F3EB", x"F48C", x"F602", x"F801", x"FA00", x"FC5A", x"FF46", x"0230", x"04C6", x"0716", x"08C3", x"0A3C", x"0BED", x"0D9E", x"0F26", x"107F", x"10F8", x"1061", x"0F57", x"0DC9", x"0B9E", x"09F3", x"08F2", x"07A1", x"0626", x"04DA", x"02DF", x"00E8", x"00B2", x"019F", x"0240", x"029B", x"01E5", x"FEF7", x"FBE3", x"FABB", x"FB10", x"FC89", x"FFBC", x"02E2", x"04A8", x"0615", x"071A", x"0694", x"0542", x"0422", x"0281", x"007A", x"FECD", x"FCEC", x"FAA7", x"F8F1", x"F7CF", x"F6E4", x"F639", x"F5A2", x"F4E4", x"F4C4", x"F510", x"F55F", x"F61E", x"F73A", x"F806", x"F92E", x"FB14", x"FC5D", x"FD49", x"FF1A", x"00F0", x"0216", x"039B", x"04EE", x"04E2", x"0574", x"07BE", x"09DE", x"0B40", x"0C11", x"0A8B", x"06B4", x"03BA", x"0278", x"021B", x"0358", x"05BA", x"06CD", x"069F", x"0617", x"0456", x"0140", x"FE7C", x"FBF9", x"F965", x"F7AF", x"F6AB", x"F59A", x"F535", x"F5D9", x"F702", x"F8FE", x"FBD3", x"FE57", x"009D", x"02C9", x"0360", x"0245", x"0085", x"FDB4", x"F9E5", x"F6C8", x"F43D", x"F102", x"EEBB", x"EE20", x"EDB5", x"ED90", x"EE78", x"EEB7", x"EE23", x"EF28", x"F1A0", x"F3DA", x"F618", x"F7AA", x"F692", x"F448", x"F36E", x"F41B", x"F656", x"FAED", x"0021", x"040E", x"074B", x"09FB", x"0B55", x"0C22", x"0D05", x"0D34", x"0CAD", x"0BF1", x"0A8F", x"08A5", x"0728", x"05DB", x"04B7", x"041C", x"0369", x"0241", x"0172", x"00D7", x"FFA3", x"FEDF", x"FED3", x"FE87", x"FEA7", x"FFC3", x"003A", x"FFA2", x"FF9B", x"FFD5", x"FFA0", x"0050", x"017F", x"0118", x"FFF4", x"FFA0", x"FEFE", x"FDD3", x"FCFF", x"FAF0", x"F6A2", x"F28D", x"F053", x"EF92", x"F0F4", x"F461", x"F728", x"F847", x"F8CC", x"F86D", x"F6E8", x"F5AC", x"F4F1", x"F3FF", x"F3A2", x"F420", x"F4CC", x"F5D7", x"F7AF", x"F9BC", x"FBF1", x"FE75", x"0091", x"0257", x"04A4", x"06E0", x"0895", x"0A70", x"0BA4", x"0B87", x"0B6F", x"0BB3", x"0B10", x"0A3B", x"0A43", x"09CD", x"08BA", x"083D", x"06F3", x"038B", x"0026", x"FDE8", x"FBAF", x"FA67", x"FA3C", x"F89B", x"F521", x"F28B", x"F150", x"F151", x"F3F9", x"F88E", x"FC74", x"FFAA", x"02CF", x"0483", x"04A4", x"0454", x"02FA", x"0075", x"FDD1", x"FB2E", x"F816", x"F58B", x"F3A7", x"F222", x"F14C", x"F0E6", x"F012", x"EFB4", x"F038", x"F0A2", x"F14E", x"F2B9", x"F390", x"F3EC", x"F574", x"F706", x"F760", x"F819", x"F947", x"F98B", x"FA3F", x"FC33", x"FCCC", x"FBD3", x"FBBF", x"FBD6", x"FB67", x"FBD6", x"FC0D", x"F936", x"F4F7", x"F1C4", x"EF4C", x"EE6B", x"F042", x"F2AD", x"F384", x"F3EB", x"F3AF", x"F20B", x"F04E", x"EF43", x"EE65", x"EE31", x"EF37", x"F055", x"F161", x"F292", x"F32F", x"F36C", x"F40B", x"F470", x"F4CE", x"F666", x"F866", x"F9AD", x"FAF4", x"FBAF", x"FA91", x"F94A", x"F8F2", x"F7EF", x"F674", x"F602", x"F54C", x"F3C7", x"F378", x"F39C", x"F206", x"F05F", x"EFEB", x"EF93", x"EFF5", x"F223", x"F347", x"F1BB", x"EF7C", x"ED7F", x"EBEC", x"ECD8", x"F085", x"F487", x"F81F", x"FBDD", x"FEE5", x"0128", x"03AC", x"05F7", x"0775", x"0882", x"08C3", x"07EE", x"06C1", x"0576", x"03F6", x"02F0", x"0223", x"0093", x"FF06", x"FDF2", x"FC86", x"FB29", x"FACD", x"FA62", x"F9C6", x"FA83", x"FBFC", x"FCAA", x"FD67", x"FE59", x"FE39", x"FE46", x"001B", x"022E", x"036E", x"0514", x"064C", x"0609", x"0594", x"04E2", x"0191", x"FBD3", x"F5F3", x"F07D", x"EC96", x"EC10", x"EDF4", x"EFD5", x"F14D", x"F26C", x"F26B", x"F1B6", x"F14C", x"F111", x"F105", x"F190", x"F276", x"F363", x"F478", x"F5C6", x"F781", x"F9F0", x"FC79", x"FEC3", x"0154", x"03FA", x"0646", x"089F", x"0AAF", x"0B0D", x"0A3B", x"094F", x"07D3", x"05F3", x"0501", x"0468", x"033E", x"02B9", x"0307", x"023C", x"0069", x"FEBD", x"FC88", x"F9F2", x"F8EF", x"F88C", x"F677", x"F355", x"F095", x"EDD7", x"EC42", x"ED54", x"EF99", x"F14F", x"F34D", x"F5D1", x"F7AE", x"F923", x"FA89", x"FAEA", x"FA08", x"F8B7", x"F6E6", x"F479", x"F204", x"F025", x"EF0F", x"EEE0", x"EF38", x"EF9C", x"F03A", x"F097", x"F0A0", x"F0CA", x"F0BA", x"EFD4", x"EEF7", x"EEA2", x"EE18", x"EDCF", x"EEA7", x"EFB7", x"F0CE", x"F357", x"F6A6", x"F8F3", x"FAFF", x"FD19", x"FE0C", x"FE90", x"0005", x"005F", x"FE2A", x"FB16", x"F81F", x"F54C", x"F4AC", x"F6F3", x"F993", x"FB57", x"FCC9", x"FD26", x"FBB6", x"F9B0", x"F78A", x"F507", x"F323", x"F292", x"F2C4", x"F377", x"F472", x"F550", x"F640", x"F75C", x"F876", x"F9F5", x"FC2B", x"FE3D", x"FFBA", x"00B5", x"FFF5", x"FD31", x"F9CD", x"F61F", x"F1C9", x"EE24", x"EBCB", x"E99B", x"E837", x"E8CF", x"E9C4", x"EA05", x"EAA2", x"EB2C", x"EAD9", x"EB95", x"EE00", x"EF70", x"EF45", x"EF02", x"EE76", x"EE61", x"F12C", x"F67F", x"FB87", x"FFF5", x"0415", x"06EE", x"0883", x"0A36", x"0BA2", x"0C35", x"0C9E", x"0D21", x"0CEB", x"0C20", x"0B1E", x"09F8", x"08F1", x"082C", x"076B", x"0698", x"0594", x"0449", x"031B", x"0245", x"0170", x"00E6", x"010A", x"0162", x"01AC", x"0270", x"02E3", x"027A", x"0234", x"0281", x"0288", x"02A9", x"036F", x"03AA", x"0349", x"03BA", x"0429", x"0285", x"FF59", x"FB96", x"F72E", x"F3E9", x"F3C7", x"F54E", x"F645", x"F6DE", x"F6C0", x"F503", x"F29D", x"F0DB", x"EF37", x"EE06", x"EE44", x"EFB5", x"F18F", x"F3F7", x"F6E1", x"F9D3", x"FD06", x"0041", x"031B", x"05C7", x"085D", x"0ABD", x"0D20", x"0F6D", x"10CE", x"1174", x"11E6", x"119D", x"10E1", x"1075", x"0F99", x"0DDB", x"0C5C", x"0B1B", x"08AA", x"05FD", x"0387", x"0050", x"FD16", x"FC04", x"FB7B", x"F9B5", x"F808", x"F6E4", x"F578", x"F5DB", x"F954", x"FD24", x"FFE3", x"0303", x"05EC", x"077B", x"08FA", x"0A70", x"0A05", x"0834", x"0682", x"0426", x"0108", x"FE1F", x"FB61", x"F89C", x"F6CB", x"F619", x"F611", x"F6DF", x"F845", x"F9A6", x"FB1F", x"FC86", x"FD60", x"FE16", x"FED7", x"FF08", x"FF36", x"FFE6", x"0042", x"00BB", x"0256", x"040C", x"0512", x"0644", x"06F0", x"0606", x"0580", x"061F", x"05CB", x"0411", x"0215", x"FEF7", x"FB4B", x"FA46", x"FBC4", x"FD6A", x"FF39", x"0127", x"016F", x"009B", x"0041", x"FFB4", x"FEBA", x"FECD", x"FFBF", x"00D9", x"0285", x"0472", x"0583", x"064E", x"0734", x"07C1", x"08DA", x"0B1E", x"0D74", x"0F7C", x"117A", x"1237", x"1176", x"1086", x"0F22", x"0CD8", x"0AEE", x"0975", x"078A", x"0647", x"0670", x"0653", x"05DB", x"05E2", x"0506", x"0351", x"0337", x"045C", x"0463", x"03A0", x"0251", x"FF6A", x"FCFE", x"FE2B", x"01A4", x"0578", x"09ED", x"0DF3", x"100C", x"117F", x"135D", x"1455", x"1469", x"1493", x"142D", x"12D2", x"1145", x"0FA0", x"0D9B", x"0C03", x"0B15", x"0A6C", x"0A2E", x"0A5B", x"0A98", x"0B0E", x"0BB9", x"0C0D", x"0C27", x"0C1E", x"0BBE", x"0BA0", x"0C58", x"0D26", x"0DE3", x"0F5F", x"10FC", x"125F", x"148B", x"16BE", x"1768", x"1718", x"16FA", x"1550", x"11AB", x"0D2D", x"0741", x"0025", x"FB25", x"F9D3", x"FA4A", x"FBD6", x"FE48", x"FF9B", x"FF46", x"FF22", x"FF2C", x"FE83", x"FE50", x"FF06", x"FFCA", x"00D9", x"02A6", x"0449", x"058C", x"071C", x"0886", x"09B0", x"0B51", x"0D2C", x"0EB1", x"1033", x"1157", x"1174", x"112D", x"10F7", x"105F", x"1007", x"104F", x"1024", x"0F8E", x"0F6D", x"0EEF", x"0D8C", x"0C50", x"0A8C", x"073B", x"042A", x"027F", x"00A3", x"FE65", x"FCC6", x"FA9B", x"F7E7", x"F789", x"F9A9", x"FC07", x"FEAC", x"01D2", x"03CE", x"04A4", x"05CF", x"0663", x"0576", x"0444", x"0339", x"01AA", x"001F", x"FEEB", x"FD70", x"FC00", x"FB3F", x"FAF2", x"FAFF", x"FB8E", x"FBDD", x"FBD8", x"FBB7", x"FB41", x"FAA1", x"FA74", x"FA83", x"FA92", x"FB67", x"FCBA", x"FDF9", x"0016", x"033D", x"064F", x"0979", x"0CFF", x"0F02", x"0F7D", x"1063", x"1154", x"1129", x"1087", x"0F0A", x"0B23", x"06DB", x"04EC", x"04B0", x"0557", x"0727", x"083B", x"06F5", x"04C5", x"028E", x"FFC2", x"FD54", x"FC55", x"FBE7", x"FBF5", x"FD67", x"FF27", x"0092", x"022A", x"038F", x"0412", x"04C2", x"05C4", x"064B", x"0654", x"0640", x"0500", x"02D8", x"007F", x"FDBB", x"FA92", x"F80F", x"F615", x"F46B", x"F3BD", x"F3BA", x"F36F", x"F355", x"F36B", x"F2C5", x"F243", x"F344", x"F4FC", x"F69F", x"F887", x"F98C", x"F907", x"F914", x"FB3A", x"FE7A", x"0255", x"06BA", x"09F3", x"0B7D", x"0CC9", x"0E28", x"0EDA", x"0F81", x"1055", x"1091", x"103B", x"1005", x"0F74", x"0E78", x"0DAE", x"0D25", x"0C81", x"0C08", x"0BB7", x"0B1A", x"0A41", x"094F", x"0824", x"06BC", x"053A", x"03D7", x"0321", x"0345", x"03E2", x"04E2", x"060B", x"069E", x"070A", x"0822", x"0922", x"0950", x"09A2", x"0A11", x"0989", x"085E", x"06E1", x"03AF", x"FF1A", x"FBEB", x"FA9F", x"FA35", x"FB07", x"FC90", x"FCA7", x"FB92", x"FAEA", x"FA09", x"F8A2", x"F81D", x"F8A9", x"F961", x"FB04", x"FD9F", x"FFB2", x"0101", x"027C", x"03D9", x"0525", x"0760", x"0A16", x"0C51", x"0E38", x"0FF2", x"10EF", x"1181", x"11F2", x"11C4", x"1101", x"100B", x"0E89", x"0CD0", x"0B41", x"0991", x"07C4", x"0662", x"04A5", x"023C", x"0073", x"FF9C", x"FEC3", x"FE49", x"FE3B", x"FD2D", x"FBD5", x"FC71", x"FEB2", x"0189", x"0544", x"090D", x"0B2D", x"0C37", x"0D19", x"0CE7", x"0B7E", x"0A20", x"086E", x"05F9", x"0394", x"0123", x"FE26", x"FB67", x"F9C1", x"F8E8", x"F933", x"FAB0", x"FC56", x"FDA2", x"FEAE", x"FF1D", x"FEF2", x"FE8F", x"FDCC", x"FC82", x"FB4C", x"FA5F", x"F9B6", x"FA36", x"FBB9", x"FD7D", x"FFB1", x"0209", x"0342", x"03AD", x"0480", x"0511", x"04C2", x"041A", x"021D", x"FDFB", x"F9D9", x"F7B8", x"F731", x"F83F", x"FAE5", x"FD04", x"FD70", x"FD6F", x"FD25", x"FC1D", x"FB4F", x"FB2E", x"FAE8", x"FAB2", x"FB81", x"FC71", x"FD3F", x"FE91", x"001B", x"014C", x"0304", x"0566", x"0756", x"08EA", x"0A43", x"0AD3", x"0A7D", x"09E1", x"08C7", x"06FD", x"051B", x"0378", x"01E6", x"0094", x"FF27", x"FD78", x"FBCD", x"FA41", x"F8B9", x"F7CA", x"F7CC", x"F811", x"F88A", x"F92B", x"F8F5", x"F7ED", x"F7BD", x"F912", x"FB97", x"FF91", x"0456", x"0859", x"0B43", x"0E02", x"101A", x"112A", x"11FE", x"123B", x"1155", x"1006", x"0EE8", x"0D44", x"0B5A", x"09F6", x"08C4", x"07D1", x"07F6", x"08F1", x"0976", x"09A9", x"0979", x"08A0", x"0750", x"066F", x"05D7", x"0595", x"064B", x"07F9", x"0A6B", x"0D4A", x"101B", x"1293", x"14AB", x"15E4", x"15E5", x"1547", x"13F0", x"11A0", x"0ECE", x"0BAD", x"072C", x"021F", x"FE65", x"FC52", x"FB87", x"FC9D", x"FE82", x"FF46", x"FF58", x"FF6F", x"FEDA", x"FDAF", x"FD72", x"FDCE", x"FE42", x"FFC7", x"01EF", x"0335", x"03D7", x"04AF", x"0567", x"0664", x"08B4", x"0B3A", x"0CDE", x"0DE6", x"0E7D", x"0E5F", x"0E21", x"0E3C", x"0E11", x"0D96", x"0D26", x"0CD2", x"0C79", x"0C20", x"0B40", x"09D9", x"07D9", x"04C4", x"0114", x"FDC8", x"FAF5", x"F899", x"F752", x"F63F", x"F44A", x"F294", x"F28F", x"F3BE", x"F639", x"FA0C", x"FD4C", x"FEA3", x"FF31", x"FF39", x"FE42", x"FD4D", x"FCE8", x"FC17", x"FB04", x"FA84", x"F9D7", x"F89A", x"F7BC", x"F71E", x"F64A", x"F61C", x"F6B1", x"F6D9", x"F67A", x"F5FD", x"F4E2", x"F37F", x"F2BC", x"F25D", x"F1FE", x"F216", x"F2D1", x"F400", x"F625", x"F906", x"FBE6", x"FE8D", x"00DF", x"0207", x"0299", x"0321", x"030E", x"021E", x"008D", x"FD8D", x"F91C", x"F50A", x"F2C3", x"F1F2", x"F2EB", x"F52B", x"F6D1", x"F73B", x"F734", x"F6B3", x"F5B0", x"F542", x"F59E", x"F637", x"F767", x"F970", x"FB47", x"FCC1", x"FE2C", x"FEF8", x"FF2F", x"FF87", x"001E", x"0031", x"000A", x"FFAC", x"FE8F", x"FCFE", x"FB6E", x"F9A9", x"F784", x"F57B", x"F3BB", x"F240", x"F11D", x"F03D", x"EF76", x"EF0A", x"EECB", x"EEDF", x"EF97", x"F0E4", x"F266", x"F46A", x"F67E", x"F7A0", x"F7D1", x"F82E", x"F8BB", x"F9D3", x"FC40", x"FF5B", x"01E0", x"042F", x"06C2", x"08BA", x"0A72", x"0C7A", x"0DF3", x"0E65", x"0EE6", x"0F39", x"0E85", x"0D73", x"0C79", x"0AD8", x"094F", x"0933", x"096A", x"08F5", x"0820", x"0695", x"03BB", x"00E2", x"FF0A", x"FD32", x"FB6A", x"FA74", x"FA0F", x"FA27", x"FB49", x"FCFB", x"FE59", x"FF57", x"0000", x"0011", x"001C", x"004E", x"0016", x"FF5E", x"FDCA", x"FA7B", x"F617", x"F227", x"EF1E", x"ED61", x"ED8F", x"EE94", x"EEDF", x"EEDD", x"EE9E", x"EDA2", x"ECAC", x"ECE5", x"EDD2", x"EF62", x"F249", x"F587", x"F7DB", x"F9C8", x"FB77", x"FC8D", x"FE26", x"0100", x"0417", x"06C6", x"0968", x"0B6C", x"0C75", x"0D51", x"0DD5", x"0D27", x"0B90", x"0965", x"06D9", x"0459", x"023F", x"003E", x"FE5C", x"FC7F", x"FA4A", x"F82F", x"F6B7", x"F589", x"F4C2", x"F4B4", x"F40E", x"F21F", x"F043", x"EF60", x"EF44", x"F0E9", x"F419", x"F68E", x"F78C", x"F836", x"F81F", x"F728", x"F6B7", x"F69D", x"F598", x"F47E", x"F3EE", x"F2D2", x"F151", x"F07E", x"EFBB", x"EED6", x"EF61", x"F10D", x"F279", x"F3C6", x"F4C5", x"F46D", x"F331", x"F271", x"F19A", x"F072", x"EFC7", x"EFA1", x"EFB1", x"F0BF", x"F2C0", x"F4D8", x"F6F1", x"F922", x"FAD5", x"FC64", x"FE14", x"FF41", x"FF8A", x"FF0B", x"FCFE", x"F986", x"F634", x"F412", x"F330", x"F43D", x"F6B8", x"F8EB", x"FA3C", x"FAFD", x"FA91", x"F905", x"F789", x"F650", x"F54F", x"F549", x"F65D", x"F792", x"F906", x"FAD1", x"FC7A", x"FE04", x"0026", x"0247", x"03CA", x"04E0", x"0559", x"04C1", x"03C7", x"02EF", x"01B5", x"0013", x"FE63", x"FC86", x"FA97", x"F90D", x"F7C1", x"F684", x"F563", x"F440", x"F30A", x"F235", x"F1C7", x"F1A2", x"F21E", x"F2F8", x"F326", x"F2E5", x"F311", x"F391", x"F4E7", x"F7DE", x"FB7C", x"FE75", x"0124", x"0376", x"0475", x"04BE", x"0506", x"0483", x"034E", x"029E", x"01CF", x"0018", x"FE6A", x"FCE0", x"FAEA", x"F9B6", x"FA50", x"FB46", x"FBF5", x"FCB2", x"FC8B", x"FB1F", x"FA27", x"FA1C", x"F9FF", x"FA39", x"FB6E", x"FCEF", x"FEF8", x"0230", x"0584", x"07BB", x"0902", x"0914", x"07E7", x"0682", x"0542", x"03B6", x"0207", x"FFD7", x"FC42", x"F813", x"F48C", x"F1FB", x"F0F5", x"F206", x"F3A1", x"F45F", x"F4A4", x"F41F", x"F245", x"F04B", x"EF27", x"EE3C", x"EE23", x"EF9C", x"F15F", x"F29A", x"F3FD", x"F524", x"F5A2", x"F6F4", x"F951", x"FB8D", x"FD9B", x"FFAD", x"00D7", x"014C", x"0245", x"034B", x"039B", x"0396", x"0324", x"01ED", x"00B1", x"FFB1", x"FE5F", x"FCC0", x"FAF7", x"F89E", x"F64D", x"F48B", x"F2F4", x"F1AF", x"F10F", x"EFBB", x"ED72", x"EB79", x"EA69", x"EA3B", x"EC4B", x"F006", x"F331", x"F568", x"F764", x"F81E", x"F7C8", x"F7D9", x"F7D0", x"F6E9", x"F67F", x"F6BD", x"F64F", x"F597", x"F545", x"F429", x"F2B9", x"F269", x"F2AF", x"F293", x"F2C8", x"F2DB", x"F1DC", x"F100", x"F128", x"F18D", x"F224", x"F36F", x"F4BF", x"F5FE", x"F823", x"FABB", x"FD29", x"FFB1", x"01FF", x"0396", x"0518", x"06B1", x"079D", x"0836", x"084C", x"068A", x"032A", x"FFA6", x"FC38", x"F998", x"F90A", x"F9D0", x"FA11", x"FA40", x"FA7B", x"F9C3", x"F8B0", x"F86C", x"F82C", x"F80B", x"F94A", x"FB63", x"FD13", x"FEE2", x"0087", x"010C", x"0140", x"020A", x"0290", x"0275", x"0254", x"016E", x"FF78", x"FDF4", x"FD0A", x"FC15", x"FB36", x"FA6D", x"F8EE", x"F74C", x"F62B", x"F53D", x"F456", x"F3D4", x"F32A", x"F272", x"F28D", x"F35A", x"F4BE", x"F724", x"F9A4", x"FAAA", x"FAB1", x"FA5F", x"F9AD", x"FA0C", x"FCA6", x"0012", x"0358", x"0731", x"0AD1", x"0D3B", x"0F88", x"11C5", x"12A5", x"12F0", x"1398", x"137A", x"1252", x"1138", x"0F7F", x"0CD1", x"0AF5", x"0A44", x"09A4", x"0961", x"0975", x"0841", x"062D", x"0497", x"033A", x"01D7", x"015E", x"0155", x"0136", x"021A", x"040C", x"0626", x"086C", x"0A8F", x"0B6E", x"0B76", x"0B74", x"0AD8", x"0A17", x"09D0", x"0870", x"051D", x"0137", x"FD4A", x"F999", x"F849", x"F96E", x"FA6E", x"FAE1", x"FB6C", x"FACC", x"F960", x"F928", x"F99E", x"F9BD", x"FAFC", x"FD7D", x"FF81", x"017E", x"0412", x"05BF", x"06D1", x"0907", x"0BB7", x"0E02", x"10A8", x"12C8", x"131C", x"12C4", x"128C", x"11C2", x"10B2", x"0FD6", x"0E26", x"0BF7", x"0A4B", x"08F8", x"07BF", x"075A", x"0703", x"0634", x"05C9", x"05A0", x"052E", x"058B", x"0696", x"0673", x"055B", x"0441", x"02B5", x"01C7", x"038B", x"06B0", x"0935", x"0BB0", x"0D98", x"0D94", x"0CED", x"0C9D", x"0B3F", x"0900", x"0792", x"0651", x"04C5", x"0471", x"04BA", x"0484", x"04B5", x"05B6", x"0656", x"06E9", x"07D4", x"07B6", x"0671", x"0530", x"03B3", x"01DC", x"00B0", x"FFB6", x"FE5B", x"FD9D", x"FDEE", x"FEA9", x"0088", x"0393", x"0630", x"084F", x"0A76", x"0B82", x"0BDC", x"0CDE", x"0D76", x"0C2D", x"09FD", x"0735", x"0373", x"0125", x"01A6", x"02E0", x"03D1", x"0503", x"053B", x"03B3", x"0290", x"01C0", x"001B", x"FECB", x"FEDD", x"FF24", x"FFC6", x"019C", x"034A", x"041C", x"055C", x"06D0", x"07BD", x"08D0", x"09C2", x"0948", x"07CE", x"0643", x"045E", x"026F", x"0134", x"FFE3", x"FE52", x"FD51", x"FCA7", x"FC0D", x"FBFA", x"FBEA", x"FB1F", x"FA50", x"F9D1", x"F944", x"F9E5", x"FC3A", x"FE90", x"0008", x"00F3", x"0084", x"FF59", x"001D", x"033C", x"06F7", x"0B3D", x"0F9F", x"122B", x"134E", x"1485", x"150E", x"1474", x"1425", x"13FC", x"1301", x"124D", x"1214", x"1135", x"1003", x"0F81", x"0EE7", x"0E44", x"0E61", x"0E60", x"0D6B", x"0C57", x"0B49", x"09FD", x"096D", x"09CE", x"0A39", x"0B03", x"0C72", x"0DBE", x"0EFC", x"109C", x"1190", x"1177", x"1130", x"101A", x"0E2D", x"0D1B", x"0CE1", x"0BD7", x"0A50", x"08A7", x"05D2", x"0361", x"03B5", x"0584", x"06E4", x"082D", x"0863", x"064A", x"0407", x"032C", x"0286", x"023C", x"0373", x"04D8", x"05A7", x"071A", x"08B9", x"0984", x"0A99", x"0C85", x"0E5B", x"1076", x"132A", x"1525", x"1623", x"1709", x"1777", x"1768", x"1792", x"1782", x"168D", x"1572", x"1418", x"121F", x"1037", x"0E7A", x"0C14", x"0990", x"0770", x"04B6", x"022A", x"0131", x"00CD", x"FFFF", x"FF6F", x"FE30", x"FB8D", x"F9E3", x"FABA", x"FC83", x"FEE9", x"023A", x"0469", x"0500", x"05A8", x"0638", x"056F", x"0473", x"03B4", x"0241", x"00F0", x"00B7", x"00A4", x"0072", x"00E2", x"0143", x"0113", x"014B", x"0199", x"0146", x"0100", x"00E4", x"0044", x"FFC0", x"FFAC", x"FF1E", x"FE6C", x"FE47", x"FE52", x"FEAD", x"0066", x"028D", x"0450", x"063D", x"078B", x"076A", x"073D", x"07EE", x"0800", x"076B", x"067F", x"03CF", x"FFBF", x"FD43", x"FCB6", x"FCBC", x"FDB0", x"FEF7", x"FE90", x"FD48", x"FCE4", x"FCB2", x"FC78", x"FD6E", x"FEF6", x"0007", x"0167", x"0305", x"03A5", x"03CD", x"041B", x"03F5", x"03BF", x"0445", x"04BC", x"0486", x"0438", x"036C", x"01D2", x"0065", x"FF45", x"FDE7", x"FCE1", x"FC8A", x"FC3B", x"FC3F", x"FCB7", x"FC99", x"FBD8", x"FB19", x"F9E4", x"F870", x"F862", x"F97D", x"FA82", x"FB74", x"FBBE", x"F9E2", x"F78A", x"F754", x"F912", x"FC4B", x"016C", x"0687", x"09D5", x"0C63", x"0EEA", x"1061", x"1146", x"1274", x"12D6", x"1229", x"11B9", x"110A", x"0FAD", x"0E89", x"0DBE", x"0C8E", x"0BA1", x"0B6A", x"0AC1", x"09BB", x"08CC", x"0751", x"056D", x"0407", x"02D0", x"017D", x"00CF", x"00C8", x"0103", x"0229", x"0400", x"0593", x"0725", x"08A4", x"08BF", x"07F3", x"0743", x"05E1", x"037C", x"0130", x"FE06", x"F989", x"F628", x"F57A", x"F60B", x"F7C3", x"FA57", x"FB3E", x"F9FA", x"F8DE", x"F826", x"F73F", x"F765", x"F8A0", x"F94D", x"F9EF", x"FB61", x"FC8A", x"FD6E", x"FF2A", x"0113", x"02AF", x"0505", x"079E", x"0952", x"0ACA", x"0C04", x"0C49", x"0C42", x"0C87", x"0C29", x"0B25", x"0A52", x"0914", x"078D", x"06B2", x"05C5", x"043F", x"02E5", x"0145", x"FE9F", x"FC68", x"FB7E", x"FAA8", x"FA2F", x"FA56", x"F908", x"F64F", x"F4EE", x"F564", x"F6D5", x"FA0D", x"FE22", x"0078", x"014E", x"0236", x"01FE", x"009C", x"FF69", x"FE17", x"FC1A", x"FB0F", x"FB32", x"FB84", x"FC4F", x"FDB6", x"FE61", x"FE6F", x"FE8E", x"FDF2", x"FC97", x"FB4E", x"F9BC", x"F794", x"F5FF", x"F4D0", x"F373", x"F2B3", x"F2C5", x"F329", x"F493", x"F762", x"FA4E", x"FD4E", x"0099", x"02C7", x"03BD", x"0500", x"0647", x"06CE", x"0787", x"078F", x"04EC", x"0126", x"FE7E", x"FCB4", x"FBFD", x"FD2A", x"FDFF", x"FCCC", x"FB27", x"F9D5", x"F844", x"F793", x"F875", x"F94D", x"F9FE", x"FB96", x"FD13", x"FE34", x"FFFA", x"01C2", x"02BD", x"03F5", x"0598", x"0682", x"0727", x"07AC", x"06C3", x"04B4", x"02F8", x"0108", x"FEEE", x"FDAD", x"FCF4", x"FC1B", x"FBEF", x"FC4A", x"FBE3", x"FB38", x"FA74", x"F8B3", x"F6D8", x"F666", x"F6B4", x"F768", x"F90D", x"F9E3", x"F87A", x"F6EB", x"F69B", x"F73E", x"F991", x"FD9F", x"00AA", x"01A7", x"0221", x"01FF", x"00FE", x"009B", x"00E8", x"007A", x"FFF9", x"FFE3", x"FF40", x"FE58", x"FDE5", x"FD23", x"FBC6", x"FAF6", x"FA5F", x"F994", x"F964", x"F9B9", x"F9B0", x"F9F2", x"FAF3", x"FBB6", x"FC88", x"FDC0", x"FEEF", x"002E", x"023C", x"0446", x"05F9", x"07E1", x"0935", x"0913", x"089A", x"07CE", x"05EA", x"0422", x"02FB", x"0074", x"FCE8", x"FA9A", x"F981", x"F964", x"FB93", x"FE72", x"FEE5", x"FDB6", x"FC41", x"F9F9", x"F7F5", x"F7E5", x"F842", x"F814", x"F899", x"F97A", x"F9C9", x"FABD", x"FC8A", x"FD7D", x"FE50", x"FFEC", x"013A", x"025C", x"045D", x"061E", x"06CA", x"07BA", x"0887", x"081A", x"071A", x"05D2", x"0341", x"0071", x"FE56", x"FC0B", x"F9CC", x"F867", x"F6BD", x"F494", x"F379", x"F2F9", x"F253", x"F28F", x"F2CF", x"F0CF", x"EDA7", x"EB8E", x"EA5F", x"EAF8", x"EE96", x"F2DC", x"F56C", x"F71E", x"F812", x"F73F", x"F5D5", x"F4B5", x"F2AF", x"F048", x"EED5", x"EDEA", x"ED8B", x"EE9A", x"F03D", x"F180", x"F2EA", x"F43C", x"F4AF", x"F53D", x"F625", x"F644", x"F638", x"F685", x"F662", x"F5F2", x"F616", x"F617", x"F5E2", x"F68B", x"F7A6", x"F887", x"FA40", x"FC79", x"FDAB", x"FEB8", x"001C", x"0084", x"00B9", x"01DE", x"01C6", x"FF42", x"FC2E", x"F933", x"F61A", x"F55A", x"F707", x"F81F", x"F7F7", x"F7B7", x"F67F", x"F4B6", x"F46F", x"F4DE", x"F48B", x"F44A", x"F434", x"F33F", x"F2CE", x"F3B7", x"F467", x"F4C4", x"F5AF", x"F606", x"F58C", x"F5A1", x"F592", x"F40D", x"F249", x"F0D4", x"EEE2", x"ED40", x"ECCF", x"EC73", x"EC25", x"ECE3", x"ED9D", x"EDE1", x"EE39", x"EE22", x"ED0C", x"EC3D", x"EC2F", x"EC34", x"ED4A", x"EF6F", x"F07C", x"F01D", x"EFB3", x"EF63", x"EFD4", x"F2EC", x"F7C3", x"FBE6", x"FF39", x"01BD", x"02AF", x"0307", x"03F6", x"04AF", x"04B9", x"04A1", x"03D2", x"021F", x"00CA", x"FFF4", x"FEE5", x"FE33", x"FDBC", x"FCA7", x"FB9C", x"FB5E", x"FB10", x"FAA1", x"FAB5", x"FAB2", x"FA19", x"F9EA", x"F9FF", x"FA24", x"FB41", x"FD30", x"FEEA", x"00AE", x"027C", x"031E", x"02E3", x"028A", x"00EB", x"FE3B", x"FC34", x"FA4B", x"F713", x"F400", x"F1C8", x"EFCE", x"EFA6", x"F295", x"F605", x"F80F", x"F967", x"F97A", x"F7FA", x"F71D", x"F794", x"F7D3", x"F81B", x"F90C", x"F980", x"F9B7", x"FB07", x"FC97", x"FD67", x"FE78", x"FF73", x"FF9C", x"0013", x"016A", x"023D", x"02D6", x"03E5", x"0496", x"0479", x"0467", x"03D7", x"026A", x"012C", x"0021", x"FEA4", x"FD47", x"FC07", x"FA44", x"F8A5", x"F7CA", x"F6D2", x"F61E", x"F671", x"F670", x"F51B", x"F3B3", x"F29A", x"F1D6", x"F33D", x"F707", x"FAD0", x"FD71", x"FF28", x"FF0E", x"FD62", x"FBBC", x"FA35", x"F857", x"F6DD", x"F5FB", x"F51E", x"F50B", x"F615", x"F74E", x"F88C", x"F9C9", x"F9DA", x"F8C9", x"F7AF", x"F63F", x"F441", x"F2C0", x"F1A5", x"F048", x"EF6B", x"EF2D", x"EEC5", x"EE9B", x"EF5A", x"F02F", x"F12C", x"F32B", x"F51E", x"F68E", x"F85F", x"F9F4", x"FA6D", x"FB53", x"FCC3", x"FCDF", x"FB95", x"F9E5", x"F72C", x"F45A", x"F410", x"F59A", x"F6FB", x"F844", x"F92E", x"F8AA", x"F7D1", x"F825", x"F870", x"F869", x"F8A7", x"F884", x"F7C1", x"F809", x"F964", x"FACA", x"FC95", x"FE68", x"FEE1", x"FE9E", x"FEB8", x"FE66", x"FD74", x"FCF7", x"FC63", x"FB3D", x"FA56", x"F9E2", x"F930", x"F902", x"F9CF", x"FAC1", x"FBAC", x"FC9D", x"FCC6", x"FC68", x"FC5F", x"FC5F", x"FC5D", x"FD3E", x"FE54", x"FE40", x"FD67", x"FC10", x"F9F1", x"F8B4", x"F9CC", x"FC31", x"FEA2", x"0122", x"02B6", x"0306", x"0347", x"0433", x"0501", x"05F1", x"0705", x"0741", x"0713", x"073D", x"0784", x"0793", x"07F4", x"07C9", x"069C", x"0575", x"04BF", x"03EE", x"0369", x"0390", x"0382", x"0334", x"034D", x"0381", x"03EA", x"0566", x"07A9", x"09FF", x"0C64", x"0E42", x"0EF4", x"0F34", x"0F57", x"0EA0", x"0DA8", x"0D5C", x"0C88", x"0ACB", x"0918", x"0736", x"0517", x"04B1", x"06A1", x"08D7", x"0A8F", x"0BE1", x"0BA7", x"0A15", x"08FE", x"0867", x"077A", x"06EA", x"06D2", x"0661", x"0632", x"0708", x"07F5", x"08E2", x"0A59", x"0BB7", x"0C9F", x"0E29", x"1010", x"117A", x"12D7", x"145A", x"150F", x"1513", x"14BB", x"135C", x"1103", x"0EBA", x"0C65", x"09F0", x"07F6", x"0627", x"0435", x"02F2", x"023E", x"015B", x"00E7", x"0124", x"0081", x"FEDD", x"FD2A", x"FB0D", x"F94B", x"FA25", x"FD5F", x"00D7", x"03EF", x"0654", x"06A4", x"05B8", x"0528", x"0479", x"033E", x"025F", x"018F", x"0074", x"004B", x"0157", x"02B6", x"0480", x"067B", x"0739", x"0700", x"06C7", x"0601", x"0496", x"03B0", x"02DE", x"01A0", x"00CD", x"0044", x"FF0E", x"FDD4", x"FD4C", x"FCF9", x"FD40", x"FEAD", x"0027", x"0136", x"0298", x"0396", x"03E8", x"0500", x"06A9", x"0747", x"071C", x"0664", x"042E", x"01E7", x"01A9", x"028F", x"0331", x"03EC", x"03EA", x"0255", x"00C2", x"001C", x"FF6F", x"FEE0", x"FEF1", x"FEAB", x"FE60", x"FF68", x"015D", x"03C5", x"06F2", x"09BB", x"0AEE", x"0B81", x"0C05", x"0BC7", x"0B82", x"0BBF", x"0B5C", x"0A5A", x"09B2", x"08FA", x"07EC", x"07D1", x"0872", x"08FA", x"09D5", x"0AA1", x"0A42", x"0978", x"08EB", x"07D8", x"06F0", x"077D", x"0841", x"0867", x"08A0", x"0839", x"0699", x"0638", x"0848", x"0B41", x"0EBC", x"12A2", x"1511", x"15D7", x"16C8", x"17D0", x"1802", x"1854", x"1881", x"178A", x"1665", x"1613", x"1592", x"14F1", x"14AD", x"1386", x"113E", x"0F63", x"0E05", x"0C6A", x"0B90", x"0B6C", x"0AD7", x"0A34", x"0A32", x"09DA", x"0962", x"09DA", x"0AE5", x"0C12", x"0DCF", x"0F38", x"0F6F", x"0F3A", x"0E8E", x"0CCD", x"0AFA", x"099D", x"0779", x"049F", x"01DA", x"FE9B", x"FB6D", x"FAB4", x"FC83", x"FF13", x"0206", x"049B", x"0534", x"0476", x"03F8", x"036B", x"02B5", x"02B7", x"0308", x"0308", x"0391", x"048F", x"0563", x"0675", x"07E0", x"08C6", x"09AE", x"0B61", x"0D28", x"0F0D", x"1186", x"13A6", x"14DE", x"15DD", x"164B", x"1575", x"143B", x"12DA", x"109C", x"0E56", x"0C94", x"0A59", x"07F4", x"064D", x"0442", x"019E", x"0019", x"FF7E", x"FE58", x"FD7C", x"FCDF", x"FB16", x"F9AA", x"FB39", x"FE8D", x"022A", x"0632", x"08F7", x"08FA", x"0828", x"07CA", x"06CD", x"0585", x"04AB", x"0319", x"00FE", x"0015", x"0025", x"0089", x"01E4", x"0320", x"02DA", x"01C4", x"00A2", x"FECC", x"FD22", x"FCA3", x"FC4E", x"FC07", x"FCB0", x"FD65", x"FD45", x"FD4A", x"FD78", x"FD58", x"FE03", x"FFEB", x"01D1", x"0406", x"06C2", x"08C5", x"0A2D", x"0C2E", x"0DF0", x"0E50", x"0DFB", x"0C5B", x"08C8", x"0588", x"0459", x"0467", x"054E", x"070A", x"07D3", x"0726", x"0643", x"0575", x"0445", x"0383", x"032C", x"02A2", x"0277", x"033D", x"0470", x"0670", x"091D", x"0AE1", x"0B78", x"0B97", x"0B14", x"0A56", x"0AAE", x"0B71", x"0B59", x"0AFD", x"0A44", x"0879", x"06AB", x"05F9", x"0572", x"0539", x"0626", x"06E0", x"06D2", x"0730", x"074E", x"062A", x"0569", x"05B3", x"05A2", x"0571", x"05BC", x"047E", x"01C9", x"0053", x"0076", x"0126", x"031F", x"05B4", x"06C8", x"06EF", x"07A7", x"082D", x"082F", x"08BE", x"0908", x"085A", x"07F4", x"07F1", x"0793", x"0750", x"0724", x"05C3", x"0382", x"0159", x"FEFF", x"FCB4", x"FB91", x"FB25", x"FAE6", x"FB87", x"FCE9", x"FE2D", x"FFE0", x"0248", x"04BC", x"0757", x"0A2C", x"0C33", x"0D25", x"0DBF", x"0D8D", x"0C91", x"0BFD", x"0BA5", x"0A74", x"08BD", x"065E", x"028F", x"FE8F", x"FCA4", x"FCD0", x"FE67", x"013A", x"03E5", x"04DA", x"0498", x"03FA", x"02B4", x"0152", x"0083", x"0023", x"0013", x"00AA", x"017F", x"025E", x"035E", x"040B", x"0413", x"03D8", x"0375", x"02EA", x"031D", x"041D", x"0512", x"05F8", x"06C5", x"0686", x"0543", x"03E9", x"0210", x"FFC7", x"FE36", x"FD64", x"FC6E", x"FC30", x"FC98", x"FBFC", x"FAC2", x"FA41", x"F9BD", x"F8B3", x"F850", x"F7A7", x"F590", x"F438", x"F56B", x"F809", x"FB6D", x"FF86", x"0214", x"0204", x"0143", x"0085", x"FF18", x"FD9B", x"FCAA", x"FB32", x"F9B1", x"F93E", x"F9A2", x"FA83", x"FC49", x"FE0A", x"FEBE", x"FED4", x"FE64", x"FD46", x"FC7D", x"FC72", x"FC74", x"FC96", x"FD1F", x"FD0B", x"FC5F", x"FBCF", x"FB26", x"FA4B", x"FA4F", x"FADB", x"FB44", x"FC28", x"FD75", x"FE2F", x"FF11", x"0101", x"02D1", x"0404", x"04DB", x"0423", x"014F", x"FEB4", x"FDA1", x"FD61", x"FE4A", x"0021", x"011A", x"009E", x"FFC5", x"FE4E", x"FBE4", x"F96E", x"F78B", x"F5F6", x"F572", x"F661", x"F842", x"FB11", x"FE44", x"00A6", x"01B2", x"018E", x"0014", x"FE3D", x"FD5F", x"FD0A", x"FCFC", x"FD6F", x"FDBC", x"FD26", x"FC99", x"FC60", x"FBBE", x"FB5B", x"FBD9", x"FC12", x"FC20", x"FCE4", x"FD68", x"FD0B", x"FD68", x"FE9C", x"FF5D", x"0044", x"0137", x"0032", x"FDD6", x"FCAF", x"FCD3", x"FDB7", x"0028", x"031F", x"0481", x"0514", x"05F2", x"0612", x"0592", x"0569", x"0525", x"0472", x"046B", x"04E3", x"050B", x"053A", x"0552", x"0485", x"034D", x"0226", x"00BA", x"FF7C", x"FF13", x"FEE6", x"FEB8", x"FF18", x"FF6C", x"FF34", x"FF4E", x"FFC6", x"003D", x"0166", x"0339", x"0476", x"0521", x"05B3", x"0527", x"03F1", x"0396", x"03AA", x"0346", x"02DB", x"0191", x"FDEA", x"F995", x"F6F8", x"F5E8", x"F670", x"F914", x"FBEC", x"FD58", x"FE4E", x"FF51", x"FF47", x"FECB", x"FE79", x"FDCD", x"FCCC", x"FC81", x"FC92", x"FCA0", x"FD14", x"FD99", x"FDA4", x"FD91", x"FD6F", x"FD29", x"FD80", x"FEC1", x"0029", x"01FE", x"0407", x"0553", x"05BE", x"05D5", x"04CC", x"02C0", x"00DB", x"FEF1", x"FCA6", x"FB1B", x"FA19", x"F833", x"F65C", x"F5B9", x"F52E", x"F4D0", x"F562", x"F532", x"F332", x"F203", x"F2F6", x"F50D", x"F8A8", x"FD5E", x"0069", x"0116", x"0158", x"0127", x"FFDF", x"FED2", x"FE1A", x"FCC7", x"FBC9", x"FBC8", x"FC18", x"FC79", x"FD42", x"FD55", x"FC5E", x"FAE0", x"F8BD", x"F656", x"F4FD", x"F48C", x"F459", x"F4CA", x"F541", x"F4AB", x"F3C9", x"F319", x"F1CC", x"F0A1", x"F0A0", x"F0D5", x"F131", x"F2CC", x"F47C", x"F514", x"F619", x"F7DB", x"F8FC", x"FA4B", x"FBF3", x"FB76", x"F8E3", x"F6FF", x"F61F", x"F5F3", x"F7D3", x"FADC", x"FC49", x"FCA2", x"FCDC", x"FBE9", x"F9BF", x"F7B2", x"F56E", x"F2A8", x"F0EB", x"F04E", x"F036", x"F10F", x"F28F", x"F388", x"F3FD", x"F3F4", x"F2F4", x"F1DB", x"F1A0", x"F1A5", x"F1EE", x"F2F7", x"F3AC", x"F3B3", x"F3E9", x"F402", x"F345", x"F2DD", x"F2F3", x"F268", x"F212", x"F273", x"F1FE", x"F0DC", x"F0C0", x"F0F7", x"F104", x"F20A", x"F2DD", x"F146", x"EEB5", x"ED2E", x"EC5A", x"ED0C", x"F048", x"F3F3", x"F650", x"F873", x"FA58", x"FB06", x"FB58", x"FBFA", x"FC26", x"FC72", x"FD9F", x"FF07", x"0045", x"0191", x"0221", x"0184", x"003C", x"FDF9", x"FAD8", x"F82D", x"F639", x"F49E", x"F415", x"F480", x"F4BA", x"F538", x"F694", x"F7BA", x"F8D9", x"FAE8", x"FCD9", x"FE20", x"FFF3", x"01C6", x"0218", x"022D", x"02D7", x"02CE", x"02B0", x"035E", x"0296", x"FF23", x"FB91", x"F90B", x"F781", x"F8A1", x"FC5C", x"FF8C", x"013C", x"02A2", x"031D", x"0253", x"01A8", x"0107", x"FF94", x"FE45", x"FDC4", x"FD72", x"FD74", x"FE15", x"FE91", x"FEB9", x"FECE", x"FE7A", x"FDF8", x"FE18", x"FEC5", x"FFB7", x"015C", x"02E6", x"03A8", x"0419", x"0431", x"0335", x"01EF", x"00D7", x"FF18", x"FD51", x"FC7F", x"FB89", x"F9DF", x"F8B4", x"F7D9", x"F68D", x"F61D", x"F68C", x"F584", x"F31B", x"F13B", x"F020", x"F01D", x"F2B2", x"F6BD", x"F9C3", x"FBE5", x"FDCB", x"FEB1", x"FEDD", x"FF22", x"FF2A", x"FE95", x"FE50", x"FE50", x"FE66", x"FEB1", x"FF2B", x"FF58", x"FF35", x"FE42", x"FC46", x"FA1B", x"F853", x"F6E8", x"F65E", x"F6A3", x"F672", x"F5D2", x"F592", x"F50E", x"F422", x"F3EB", x"F3C8", x"F2F9", x"F2DC", x"F3F4", x"F4AF", x"F562", x"F708", x"F83E", x"F8F2", x"FAA5", x"FC19", x"FAFA", x"F865", x"F5C1", x"F2DF", x"F133", x"F264", x"F471", x"F564", x"F60E", x"F62E", x"F4E1", x"F310", x"F1C0", x"F043", x"EF15", x"EF56", x"F096", x"F245", x"F48C", x"F6F1", x"F8D5", x"FA45", x"FAFB", x"FAD5", x"FA71", x"FA49", x"FA88", x"FB9A", x"FD40", x"FE8F", x"FF78", x"0001", x"FFA2", x"FECC", x"FE3A", x"FD6E", x"FC58", x"FBF5", x"FBE0", x"FB4B", x"FB0A", x"FB83", x"FBC1", x"FC75", x"FE60", x"FFAA", x"FF22", x"FE09", x"FCF5", x"FBE9", x"FC8F", x"FF43", x"01F9", x"03B7", x"0555", x"065C", x"067D", x"069A", x"0711", x"0734", x"078C", x"0865", x"093D", x"0996", x"098A", x"0920", x"085B", x"0747", x"05B7", x"03D3", x"01EF", x"0021", x"FF12", x"FF13", x"FF60", x"FFAA", x"0048", x"00D7", x"011A", x"01D9", x"0312", x"0386", x"03D8", x"04BD", x"051C", x"04CF", x"0501", x"050D", x"0431", x"03CE", x"03EC", x"020F", x"FE1A", x"F9D6", x"F584", x"F21B", x"F225", x"F4E3", x"F795", x"F9CD", x"FC0E", x"FD09", x"FCEB", x"FCF0", x"FC9B", x"FB61", x"FA8B", x"FAD4", x"FB80", x"FCB8", x"FEAB", x"0095", x"0223", x"0372", x"0435", x"0452", x"0465", x"04B9", x"05A9", x"0756", x"0935", x"0AAB", x"0B9C", x"0B76", x"0A06", x"0808", x"057E", x"023F", x"FF44", x"FD48", x"FB51", x"F995", x"F8BE", x"F7F2", x"F704", x"F763", x"F87D", x"F848", x"F73E", x"F683", x"F5CE", x"F61F", x"F911", x"FD0E", x"FFCE", x"01C4", x"031C", x"0300", x"0203", x"0161", x"008A", x"FF72", x"FF40", x"FFE1", x"0053", x"00A0", x"00D1", x"00A8", x"0025", x"FF78", x"FE6C", x"FD2E", x"FC07", x"FB4D", x"FB63", x"FC05", x"FC69", x"FCBC", x"FD0D", x"FCE6", x"FCD9", x"FD7A", x"FDF7", x"FE0C", x"FEF3", x"0032", x"00E3", x"01C2", x"0313", x"036B", x"03D5", x"05A5", x"0724", x"06C8", x"05B3", x"041A", x"01BA", x"0116", x"035B", x"0623", x"0838", x"0A5A", x"0B62", x"0A9F", x"098C", x"085B", x"0614", x"03AF", x"026C", x"018C", x"0117", x"0199", x"026A", x"0321", x"0427", x"0501", x"0522", x"04FB", x"04A5", x"043A", x"0465", x"0559", x"0646", x"0752", x"082D", x"080C", x"0746", x"0689", x"0549", x"03CD", x"033A", x"02C0", x"01C8", x"0152", x"0127", x"005F", x"0049", x"0172", x"0192", x"FFFF", x"FE12", x"FB90", x"F906", x"F91F", x"FBAB", x"FE10", x"FFD9", x"018C", x"01F0", x"0151", x"015D", x"01AF", x"0190", x"0211", x"0383", x"04AB", x"0576", x"05E0", x"0552", x"03DB", x"021D", x"0009", x"FDD4", x"FC03", x"FAE4", x"FADE", x"FC51", x"FE99", x"0145", x"044E", x"06E1", x"08C8", x"0AD7", x"0CA6", x"0D99", x"0EC4", x"106C", x"115C", x"11F1", x"12C2", x"1257", x"10C3", x"103F", x"1034", x"0EB8", x"0C90", x"0A2B", x"06AD", x"0430", x"0560", x"087D", x"0B6F", x"0E9D", x"111A", x"1193", x"119E", x"121E", x"118D", x"1005", x"0EDF", x"0D9E", x"0C23", x"0B61", x"0B06", x"0A38", x"098B", x"08E9", x"07AD", x"0671", x"0587", x"04C2", x"04AD", x"05AF", x"06DB", x"0830", x"09CF", x"0AA4", x"0A84", x"0A33", x"08EB", x"0693", x"04C9", x"03C1", x"028D", x"0226", x"02A5", x"0232", x"01B3", x"02B6", x"03B0", x"02FE", x"01B5", x"FF77", x"FBB7", x"F990", x"FABB", x"FD29", x"FFB5", x"02E4", x"0511", x"0578", x"05D3", x"0652", x"05D6", x"0543", x"0589", x"05D4", x"05F7", x"0647", x"0636", x"057E", x"049B", x"0354", x"018E", x"FFA6", x"FDCE", x"FC86", x"FC83", x"FD51", x"FE4F", x"FFA8", x"009C", x"008E", x"0067", x"0059", x"FF5D", x"FE71", x"FEC6", x"FF54", x"0010", x"020C", x"03A8", x"03B4", x"0432", x"05CC", x"0672", x"0654", x"05FD", x"03B9", x"004A", x"FF2E", x"0053", x"01B8", x"037E", x"051D", x"048B", x"02B2", x"0179", x"000D", x"FE51", x"FD87", x"FD61", x"FD20", x"FD52", x"FDE2", x"FDF8", x"FE24", x"FE71", x"FE32", x"FD97", x"FCD8", x"FB9C", x"FA86", x"FA62", x"FA87", x"FAEF", x"FC1A", x"FD1A", x"FD8D", x"FE81", x"FF7A", x"FF89", x"FFE8", x"00DB", x"0118", x"0140", x"022E", x"0230", x"0161", x"0204", x"038A", x"040D", x"0436", x"0386", x"007D", x"FD1D", x"FC5E", x"FD5F", x"FEED", x"0179", x"03CF", x"047D", x"04EF", x"061D", x"06DE", x"0779", x"08AB", x"09E1", x"0AAC", x"0B73", x"0BDA", x"0B8E", x"0AF9", x"09EC", x"0850", x"0655", x"0411", x"01DA", x"00AC", x"0089", x"00EB", x"0219", x"03A0", x"047A", x"054A", x"067A", x"06F2", x"06DD", x"0783", x"0850", x"08DA", x"0A96", x"0C93", x"0CE9", x"0C90", x"0CD6", x"0C55", x"0AD6", x"097E", x"06E4", x"02C2", x"003E", x"00F7", x"0358", x"0701", x"0B61", x"0E15", x"0E83", x"0E79", x"0DFF", x"0CA7", x"0B7A", x"0B01", x"0A8A", x"0A66", x"0AD7", x"0B24", x"0B53", x"0B9D", x"0BA5", x"0B53", x"0AEB", x"0A3F", x"09B3", x"0A11", x"0AEF", x"0C08", x"0D88", x"0E97", x"0E83", x"0E20", x"0D4D", x"0B38", x"08A6", x"068F", x"0416", x"01CD", x"00E5", x"FFFC", x"FE05", x"FCD7", x"FCE2", x"FCF0", x"FD61", x"FE70", x"FDCC", x"FBC8", x"FB34", x"FC92", x"FE9D", x"01CA", x"0550", x"06EA", x"0703", x"0711", x"06A9", x"0598", x"0510", x"04F5", x"0483", x"03F7", x"0359", x"0234", x"00B0", x"FF65", x"FDFF", x"FC66", x"FAA3", x"F89C", x"F6FE", x"F63D", x"F63E", x"F6FE", x"F83A", x"F8D5", x"F8BA", x"F880", x"F7BF", x"F655", x"F56D", x"F53E", x"F513", x"F606", x"F84E", x"FA11", x"FB1F", x"FD09", x"FF34", x"00A4", x"0230", x"02FC", x"012A", x"FE6C", x"FD80", x"FE10", x"FF9F", x"0282", x"04FC", x"0511", x"03E7", x"025B", x"FFDC", x"FCF4", x"FAEF", x"F973", x"F850", x"F7E2", x"F7E0", x"F7AE", x"F79C", x"F7C6", x"F7E3", x"F7F8", x"F7D6", x"F7A9", x"F80E", x"F94E", x"FB17", x"FD82", x"FFD1", x"00E0", x"0133", x"0141", x"0070", x"FF0D", x"FE19", x"FCD0", x"FAE5", x"F9DE", x"F95E", x"F7E1", x"F67B", x"F686", x"F6B0", x"F6EE", x"F815", x"F832", x"F5EE", x"F3F7", x"F3E7", x"F4F1", x"F767", x"FB62", x"FE64", x"FFA9", x"00DC", x"0239", x"0301", x"0433", x"0619", x"0787", x"086A", x"091A", x"08B8", x"0736", x"054C", x"030E", x"00A2", x"FE7C", x"FCB2", x"FB5F", x"FB24", x"FC01", x"FDCA", x"0085", x"039D", x"0633", x"08BA", x"0AF0", x"0C17", x"0CBD", x"0D5C", x"0D60", x"0D28", x"0DE2", x"0E5E", x"0DA7", x"0CF1", x"0C9F", x"0B85", x"0A61", x"0962", x"06BD", x"028D", x"FFCB", x"FF48", x"0084", x"03EE", x"089E", x"0C0E", x"0DE8", x"0F5B", x"0FE2", x"0F3F", x"0E8F", x"0E1A", x"0D4E", x"0C83", x"0BD0", x"0AA5", x"0909", x"0794", x"065F", x"0555", x"0453", x"0321", x"0218", x"017D", x"0197", x"02AD", x"0495", x"0625", x"0736", x"07EB", x"07A6", x"0637", x"04AE", x"030A", x"00DA", x"FF81", x"FF6C", x"FEC9", x"FD69", x"FC9D", x"FBC2", x"FA86", x"FA51", x"FA60", x"F862", x"F59C", x"F467", x"F4BB", x"F69E", x"FB10", x"FFF7", x"02E7", x"04C9", x"065B", x"06C3", x"0686", x"06D7", x"06BF", x"05C4", x"04D5", x"039A", x"0158", x"FEE5", x"FC7E", x"F9C0", x"F6E7", x"F46B", x"F1DD", x"EFBC", x"EEAE", x"EE8C", x"EF3B", x"F0AB", x"F1D2", x"F24C", x"F26F", x"F1F3", x"F10F", x"F0E0", x"F161", x"F1F7", x"F363", x"F54A", x"F5D8", x"F57E", x"F581", x"F549", x"F4A8", x"F4D5", x"F43B", x"F13B", x"EDDA", x"EC26", x"EBAF", x"ECE4", x"F054", x"F35B", x"F48B", x"F51B", x"F56B", x"F4AB", x"F413", x"F482", x"F52C", x"F61D", x"F7DC", x"F986", x"FA94", x"FB9A", x"FC73", x"FD06", x"FD63", x"FD65", x"FD0B", x"FCF1", x"FD56", x"FE3C", x"FFEE", x"01B9", x"02E9", x"042E", x"0591", x"0652", x"06F5", x"07DF", x"079B", x"06BD", x"06B1", x"0679", x"0517", x"0456", x"045F", x"03F2", x"0461", x"05DF", x"0565", x"0263", x"FF9B", x"FD79", x"FC43", x"FDDC", x"017B", x"03DC", x"050C", x"0622", x"0634", x"05A1", x"0620", x"06F1", x"0753", x"082B", x"0925", x"0918", x"0886", x"07B7", x"05EC", x"03D1", x"01F3", x"FFEB", x"FDDC", x"FCA3", x"FBB2", x"FB13", x"FB77", x"FC33", x"FCBD", x"FD99", x"FE41", x"FDDF", x"FD6A", x"FD28", x"FC78", x"FC4C", x"FD85", x"FE4F", x"FE43", x"FE7C", x"FE41", x"FCFE", x"FC17", x"FB10", x"F7D1", x"F365", x"F01C", x"EE22", x"EE15", x"F0F4", x"F4E7", x"F77F", x"F920", x"FA2A", x"FA25", x"F9F7", x"FAB0", x"FBD9", x"FD21", x"FEAC", x"FFD1", x"001A", x"FFF4", x"FFAC", x"FF6E", x"FF7A", x"FF4F", x"FEB7", x"FE01", x"FD43", x"FCA9", x"FCDB", x"FD8A", x"FDD2", x"FE03", x"FE34", x"FD68", x"FC08", x"FAE8", x"F911", x"F6AC", x"F56D", x"F4DF", x"F3A4", x"F2AA", x"F28D", x"F22C", x"F28B", x"F4E3", x"F6E6", x"F687", x"F535", x"F39B", x"F1C0", x"F1B9", x"F439", x"F6B1", x"F7DB", x"F8BA", x"F8C8", x"F7EA", x"F7AF", x"F829", x"F821", x"F7E4", x"F7DB", x"F716", x"F5E9", x"F50E", x"F40A", x"F2A0", x"F16A", x"F006", x"EE54", x"ED44", x"ED1A", x"ED95", x"EF11", x"F11D", x"F287", x"F357", x"F38E", x"F2BA", x"F1A0", x"F13E", x"F12F", x"F1B2", x"F3BB", x"F65F", x"F841", x"FA45", x"FC5C", x"FD86", x"FECB", x"00A0", x"00DB", x"FEBD", x"FC3E", x"FA01", x"F871", x"F968", x"FC7F", x"FF27", x"0092", x"014B", x"009B", x"FEDA", x"FD94", x"FCF1", x"FC95", x"FCE8", x"FD8E", x"FD8F", x"FCFF", x"FC1D", x"FAE5", x"F9E4", x"F96A", x"F92D", x"F9B4", x"FB37", x"FD57", x"FFFD", x"02F8", x"04F3", x"05C1", x"0628", x"05EB", x"04FF", x"0481", x"03DA", x"01E2", x"FFCB", x"FE4A", x"FBF7", x"F95F", x"F7DD", x"F686", x"F54F", x"F625", x"F800", x"F817", x"F6F3", x"F588", x"F38B", x"F28C", x"F4A1", x"F801", x"FAAA", x"FCEE", x"FE63", x"FE41", x"FDFE", x"FE86", x"FF05", x"FFA4", x"00A9", x"0105", x"005C", x"FF61", x"FDFF", x"FC2E", x"FAF7", x"FA0A", x"F909", x"F879", x"F877", x"F8A8", x"F99D", x"FB91", x"FD94", x"FFB4", x"0200", x"0371", x"03FF", x"045D", x"040A", x"0311", x"02D6", x"0364", x"0395", x"0409", x"04DE", x"04E8", x"048D", x"04D5", x"0458", x"01ED", x"FEEE", x"FC56", x"FAAD", x"FB93", x"FFA3", x"049F", x"08DB", x"0BF2", x"0D4D", x"0CAF", x"0B6A", x"0A30", x"08F9", x"07ED", x"06E9", x"053B", x"02E8", x"0042", x"FDCC", x"FBFD", x"FAFB", x"FA3E", x"F998", x"F921", x"F8BA", x"F8E9", x"F9F8", x"FB6E", x"FCAC", x"FDCF", x"FE4F", x"FDD1", x"FD30", x"FC84", x"FB46", x"FA02", x"F985", x"F8FA", x"F7FD", x"F75C", x"F6C7", x"F5C4", x"F5A3", x"F6E2", x"F79C", x"F715", x"F632", x"F4FF", x"F40B", x"F553", x"F8EA", x"FCBF", x"003F", x"0364", x"0560", x"0642", x"0712", x"07D5", x"07D7", x"07B0", x"073A", x"0603", x"0443", x"02AD", x"00F1", x"FF3A", x"FDAC", x"FBD4", x"F980", x"F763", x"F5B8", x"F4B6", x"F4CE", x"F592", x"F65B", x"F70B", x"F789", x"F799", x"F803", x"F906", x"FA1E", x"FB99", x"FDD0", x"FFA4", x"00AC", x"0197", x"01F3", x"0141", x"00E0", x"00BA", x"FED7", x"FB54", x"F7BA", x"F41F", x"F19D", x"F223", x"F4E5", x"F789", x"F9D8", x"FBC1", x"FC28", x"FBAA", x"FBBB", x"FC10", x"FC94", x"FDFD", x"FFA4", x"005E", x"0048", x"FF82", x"FDD9", x"FC25", x"FB14", x"FA48", x"FA0F", x"FAA8", x"FBB2", x"FD23", x"FF2C", x"0119", x"02A3", x"0418", x"051A", x"0597", x"0648", x"06B9", x"0641", x"05C0", x"0539", x"03B1", x"01D3", x"00A8", x"FF68", x"FE91", x"FF8C", x"00DA", x"0068", x"FED5", x"FCC0", x"FA1E", x"F8D0", x"FA82", x"FD6F", x"0023", x"02E8", x"050B", x"05F8", x"06DF", x"0876", x"0A14", x"0BED", x"0E2D", x"0F95", x"0FAB", x"0EBE", x"0CB5", x"0A03", x"0787", x"0537", x"02CA", x"00BF", x"FEFF", x"FD69", x"FCE0", x"FD5A", x"FE55", x"FFF8", x"01F8", x"0355", x"040C", x"04B2", x"048F", x"0410", x"04AC", x"05E1", x"06CD", x"0817", x"097F", x"09B1", x"0998", x"0A15", x"093E", x"062A", x"028C", x"FEE0", x"FBD1", x"FBBE", x"FEFD", x"02F6", x"0648", x"0921", x"0A60", x"0A2D", x"0A2F", x"0AB7", x"0B12", x"0BC2", x"0CA3", x"0CA3", x"0BCD", x"0ACC", x"0960", x"0804", x"073F", x"06B3", x"05FA", x"057E", x"0520", x"04A8", x"04C6", x"0563", x"05EE", x"067A", x"06D2", x"0639", x"050C", x"03B1", x"01CC", x"FFD1", x"FEBC", x"FDD5", x"FCC6", x"FC84", x"FCF3", x"FD8E", x"FF9E", x"031C", x"05A5", x"065A", x"062E", x"04D0", x"030F", x"034A", x"0569", x"0774", x"0965", x"0B6F", x"0C61", x"0C8F", x"0D0D", x"0D52", x"0CD2", x"0C6F", x"0BDD", x"0A7A", x"08F7", x"07A1", x"05FF", x"04A2", x"0393", x"020C", x"003F", x"FEC4", x"FD47", x"FC30", x"FC30", x"FCA2", x"FD00", x"FDC1", x"FE24", x"FDB0", x"FD5C", x"FD3E", x"FCBB", x"FD3B", x"FF41", x"014E", x"0353", x"05F0", x"0784", x"07E2", x"0918", x"0A26", x"08E0", x"0632", x"0303", x"FEA2", x"FB71", x"FBE2", x"FE04", x"FFE3", x"0206", x"0333", x"023E", x"012C", x"00E0", x"0039", x"FFE3", x"0096", x"00E8", x"0069", x"001D", x"FF18", x"FD3A", x"FC06", x"FBA3", x"FB88", x"FCC2", x"FF07", x"00F1", x"02A0", x"0456", x"04EF", x"04E5", x"04EF", x"0443", x"02F6", x"0223", x"0114", x"FF8D", x"FEE3", x"FE9C", x"FD65", x"FC41", x"FB7A", x"F9EB", x"F913", x"FA92", x"FC37", x"FC9B", x"FC79", x"FB36", x"F8A9", x"F7DD", x"F9DD", x"FC82", x"FF51", x"024B", x"03F5", x"0469", x"0570", x"06D4", x"080E", x"09C5", x"0B81", x"0C28", x"0C3E", x"0BF3", x"0B00", x"0A24", x"09D7", x"0939", x"0876", x"0800", x"0743", x"06A5", x"0735", x"0847", x"0999", x"0BBB", x"0DE7", x"0F28", x"104C", x"1116", x"1049", x"0F31", x"0F1D", x"0F0C", x"0F29", x"1086", x"1146", x"105E", x"0FE4", x"1000", x"0E98", x"0C35", x"09BC", x"062F", x"0333", x"0411", x"0815", x"0CE6", x"11FE", x"1616", x"1743", x"16C5", x"1641", x"154B", x"13ED", x"1302", x"11AC", x"0F48", x"0CBD", x"0A15", x"0726", x"04BB", x"032C", x"01C0", x"00C8", x"0093", x"0085", x"00E1", x"020F", x"037E", x"04CC", x"064C", x"0739", x"0757", x"0749", x"06D5", x"057A", x"0443", x"03A0", x"02AB", x"01F8", x"0208", x"01A0", x"00E1", x"019F", x"0353", x"0430", x"0488", x"044F", x"0273", x"00C0", x"0175", x"03C2", x"065A", x"09A8", x"0CD8", x"0EB3", x"1009", x"1176", x"11F2", x"11AB", x"114B", x"1059", x"0E91", x"0C96", x"0A5C", x"07F1", x"060B", x"0487", x"02DE", x"0140", x"FF77", x"FD7B", x"FC13", x"FBA5", x"FBB1", x"FC72", x"FDC2", x"FEAA", x"FF52", x"004F", x"0080", x"FFDF", x"FFDD", x"0018", x"FFE2", x"0065", x"012B", x"0048", x"FEF2", x"FEEA", x"FE95", x"FD0C", x"FB7A", x"F8D8", x"F49C", x"F224", x"F2E2", x"F4C2", x"F718", x"FA08", x"FB62", x"FAF9", x"FB14", x"FBAF", x"FBF3", x"FCED", x"FE81", x"FF21", x"FF2B", x"FF08", x"FDC1", x"FBDA", x"FAA1", x"F9CF", x"F981", x"FAB2", x"FCB2", x"FEAC", x"013B", x"040D", x"064B", x"0895", x"0ADE", x"0C25", x"0CFC", x"0DCD", x"0DAE", x"0D1A", x"0D2C", x"0CDD", x"0BCC", x"0B10", x"09E4", x"078E", x"064E", x"06EE", x"077D", x"077D", x"071D", x"04B8", x"00E2", x"FEEB", x"FF30", x"0041", x"0252", x"04D4", x"0625", x"06F0", x"08A9", x"0AB9", x"0CD6", x"0F84", x"11FC", x"133C", x"13A7", x"1317", x"115F", x"0F4F", x"0D34", x"0AAE", x"0804", x"0569", x"0289", x"0011", x"FEA9", x"FDE2", x"FDCC", x"FE78", x"FEF6", x"FF08", x"FF60", x"FF57", x"FE70", x"FDF0", x"FE23", x"FE51", x"FF85", x"01D7", x"0320", x"0317", x"036F", x"037E", x"0232", x"00A2", x"FE92", x"FAAE", x"F743", x"F713", x"F929", x"FC54", x"00AA", x"0439", x"055C", x"05BA", x"0669", x"067B", x"0666", x"0705", x"0721", x"0655", x"05B3", x"04BF", x"02E2", x"0121", x"FFE6", x"FE8D", x"FDA6", x"FD96", x"FD66", x"FCF1", x"FD08", x"FD34", x"FD5F", x"FDD9", x"FE4D", x"FE24", x"FDF4", x"FD90", x"FC96", x"FBC9", x"FB49", x"FA7E", x"FA35", x"FAAA", x"FA98", x"FA8B", x"FBF3", x"FDAC", x"FE5C", x"FE83", x"FD30", x"F948", x"F590", x"F47E", x"F4E8", x"F67A", x"F9F7", x"FD61", x"FF81", x"01FB", x"049E", x"059A", x"05AC", x"05BE", x"04A9", x"02E3", x"01D3", x"006C", x"FE5E", x"FCDA", x"FBC0", x"FA4A", x"F92A", x"F845", x"F6A6", x"F528", x"F49A", x"F498", x"F570", x"F725", x"F871", x"F956", x"FA33", x"FA4E", x"FA15", x"FB03", x"FC74", x"FE0F", x"0102", x"03D8", x"048B", x"050E", x"0671", x"06AA", x"060E", x"0591", x"02AE", x"FD9C", x"FAF0", x"FB3B", x"FC76", x"FF5B", x"02F8", x"03CF", x"02D5", x"02F9", x"02DE", x"0209", x"0266", x"02C0", x"0183", x"0073", x"FFD4", x"FDE1", x"FBBD", x"FAC8", x"F9F4", x"F9E2", x"FBF5", x"FE87", x"00A0", x"02FA", x"04B9", x"0525", x"0593", x"05CD", x"04F6", x"0421", x"035D", x"0155", x"FF2F", x"FDBE", x"FB83", x"F918", x"F799", x"F506", x"F11E", x"EEFB", x"EE85", x"EE1B", x"EECB", x"EFA6", x"ED90", x"EA2C", x"E923", x"E98E", x"EAF4", x"EE8B", x"F236", x"F3B5", x"F520", x"F75D", x"F8DF", x"FA2B", x"FC1B", x"FD02", x"FCEB", x"FD51", x"FDA2", x"FD48", x"FD66", x"FD7A", x"FCA1", x"FBCC", x"FB08", x"F9C3", x"F901", x"F940", x"F9AF", x"FAB9", x"FC9C", x"FE01", x"FF0C", x"0072", x"00CA", x"FFD9", x"FF3E", x"FEC8", x"FE10", x"FF2F", x"01AB", x"02C4", x"033B", x"0466", x"04AA", x"03EC", x"03FA", x"02EE", x"FF66", x"FCDA", x"FD22", x"FED2", x"0232", x"0734", x"0A34", x"0A43", x"09CB", x"08CC", x"06B8", x"0567", x"04FC", x"03C1", x"0275", x"01CD", x"0055", x"FE0B", x"FC1F", x"F9F5", x"F774", x"F60E", x"F576", x"F4DD", x"F4E8", x"F591", x"F5DB", x"F672", x"F781", x"F80C", x"F858", x"F8E8", x"F8AA", x"F7CC", x"F77A", x"F6E2", x"F5EC", x"F5F0", x"F60F", x"F4C7", x"F3FC", x"F4B7", x"F56E", x"F691", x"F878", x"F827", x"F503", x"F273", x"F164", x"F134", x"F37D", x"F7CB", x"FAE8", x"FD1D", x"001A", x"0265", x"0397", x"0517", x"05F3", x"04FE", x"03EB", x"0309", x"011D", x"FF0B", x"FD76", x"FB1B", x"F870", x"F682", x"F45E", x"F1D3", x"F02B", x"EEFB", x"EE1E", x"EEEE", x"F0DD", x"F2D9", x"F552", x"F7BD", x"F880", x"F8C0", x"F92C", x"F8C0", x"F87D", x"F996", x"F9C6", x"F853", x"F782", x"F6C6", x"F4F2", x"F3ED", x"F312", x"EF3E", x"EA4F", x"E782", x"E63C", x"E6BE", x"EA8B", x"EEA5", x"F049", x"F169", x"F2E3", x"F370", x"F499", x"F71A", x"F87F", x"F892", x"F8CB", x"F810", x"F5FB", x"F452", x"F2A1", x"F021", x"EEA5", x"EE8E", x"EEE8", x"F070", x"F358", x"F5D2", x"F808", x"FA87", x"FC3A", x"FD35", x"FED1", x"FFC8", x"FFA4", x"FFA3", x"FF0A", x"FD0F", x"FB94", x"FA97", x"F804", x"F51F", x"F383", x"F1CC", x"F093", x"F169", x"F1AD", x"EF44", x"ECAC", x"EB0B", x"E9DE", x"EB1F", x"EF44", x"F30A", x"F598", x"F898", x"FB37", x"FD1D", x"FFD7", x"02A2", x"03A5", x"03C5", x"038D", x"020B", x"0026", x"FEC8", x"FCF9", x"FAB5", x"F905", x"F780", x"F5DD", x"F534", x"F534", x"F55A", x"F632", x"F77D", x"F83C", x"F8ED", x"F98F", x"F960", x"F8FE", x"F91C", x"F904", x"F942", x"FB3D", x"FD9C", x"FF3D", x"00EA", x"022F", x"01E7", x"0189", x"01A6", x"003E", x"FD3F", x"FB30", x"FA31", x"FA8B", x"FDCB", x"02D5", x"06AB", x"090F", x"0AC6", x"0AFF", x"0A46", x"0A33", x"0A2A", x"0965", x"08E1", x"0893", x"076F", x"0610", x"04E8", x"0346", x"019B", x"00C4", x"003C", x"FFA2", x"FF73", x"FF46", x"FEC3", x"FE85", x"FE5B", x"FDD8", x"FD63", x"FCFD", x"FC39", x"FBB3", x"FB90", x"FB0C", x"FADA", x"FBB8", x"FC55", x"FC59", x"FD0D", x"FDD0", x"FDF0", x"FEC8", x"FFA7", x"FDC8", x"F9C0", x"F61D", x"F2B4", x"F0AB", x"F20C", x"F522", x"F72B", x"F93A", x"FBB7", x"FD1E", x"FE0C", x"FF95", x"FFD7", x"FE91", x"FDBC", x"FD28", x"FBF0", x"FB65", x"FB2E", x"F9CF", x"F80E", x"F6BE", x"F4CF", x"F2A1", x"F159", x"F058", x"EFAE", x"F072", x"F207", x"F390", x"F58E", x"F77D", x"F895", x"F9D6", x"FB4B", x"FC41", x"FDC1", x"0036", x"01BE", x"0294", x"03A9", x"03D0", x"02EC", x"02B4", x"01AF", x"FDF7", x"F9B6", x"F695", x"F44D", x"F45F", x"F7AC", x"FB02", x"FCA2", x"FDFA", x"FE90", x"FE0B", x"FE2B", x"FF10", x"FEED", x"FE59", x"FDFD", x"FCB5", x"FAF3", x"F9C0", x"F851", x"F666", x"F557", x"F4AD", x"F40F", x"F485", x"F5BD", x"F696", x"F7C6", x"F950", x"FA51", x"FB7B", x"FD7D", x"FEE0", x"FFC0", x"009E", x"0039", x"FE7C", x"FD3C", x"FBD8", x"F919", x"F6A5", x"F4E2", x"F2A3", x"F17D", x"F277", x"F2BE", x"F148", x"F006", x"EEF3", x"EDF4", x"EF99", x"F3A5", x"F715", x"F9FE", x"FD37", x"FF89", x"010B", x"0368", x"0587", x"065E", x"074A", x"0864", x"089B", x"08CB", x"0956", x"08BF", x"0773", x"0671", x"0532", x"03C3", x"0371", x"03D6", x"0458", x"05F3", x"0873", x"0AC8", x"0D09", x"0F1A", x"0FD5", x"0F7D", x"0EE5", x"0DA9", x"0C54", x"0C33", x"0C88", x"0C9D", x"0D3F", x"0DF5", x"0DCD", x"0DF2", x"0E8B", x"0DDB", x"0C35", x"0B7B", x"0B84", x"0CA7", x"101D", x"1483", x"174E", x"18CE", x"197E", x"188B", x"1705", x"161C", x"14DE", x"1306", x"1185", x"0FC9", x"0D27", x"0ABC", x"0849", x"0533", x"0273", x"00BF", x"FF4C", x"FECF", x"FFCE", x"0100", x"020B", x"03B6", x"052F", x"05E7", x"0712", x"0822", x"083F", x"0878", x"08F9", x"08A0", x"0881", x"093F", x"0918", x"0833", x"0828", x"0804", x"07A9", x"08F3", x"0A6A", x"093F", x"06B6", x"0436", x"0101", x"FF3D", x"00CE", x"0328", x"0499", x"06BE", x"08D7", x"09C1", x"0B52", x"0D71", x"0DAD", x"0CD5", x"0C42", x"0AB9", x"08C5", x"0812", x"0701", x"0488", x"0255", x"0023", x"FCFA", x"FABC", x"F9AB", x"F813", x"F6CB", x"F6FD", x"F73E", x"F7B5", x"F957", x"FA8F", x"FA6E", x"FA59", x"F9DF", x"F88C", x"F833", x"F8E9", x"F8F9", x"F923", x"F9E1", x"F97A", x"F8BC", x"F8EB", x"F7F5", x"F4E1", x"F1C6", x"EEE7", x"EC5D", x"ECD4", x"F052", x"F401", x"F787", x"FB39", x"FD83", x"FED8", x"00FB", x"02D4", x"03AD", x"04BF", x"0578", x"04F1", x"04A3", x"049C", x"038A", x"026D", x"0212", x"0180", x"01AD", x"03F5", x"06E2", x"098C", x"0CC0", x"0F5F", x"10A1", x"1260", x"14B3", x"1635", x"17C0", x"1955", x"1926", x"181F", x"17D9", x"16FA", x"1528", x"13FD", x"1248", x"0F47", x"0D55", x"0C8B", x"0A6E", x"078A", x"0526", x"0228", x"FFEC", x"011C", x"044E", x"0764", x"0B12", x"0ED5", x"1116", x"133E", x"15FD", x"1785", x"17DE", x"1805", x"171D", x"1514", x"136C", x"11AB", x"0EDA", x"0C15", x"0962", x"05F2", x"02C7", x"00B5", x"FEAD", x"FCF1", x"FC6B", x"FC3B", x"FC2D", x"FD14", x"FE43", x"FEC2", x"FF63", x"FFE3", x"FFA2", x"FFB3", x"00D6", x"01CA", x"02DB", x"0489", x"0597", x"05E6", x"06D5", x"07A3", x"06C3", x"0566", x"0440", x"030C", x"035B", x"065B", x"0A2C", x"0D57", x"103D", x"11FB", x"1216", x"11C2", x"1156", x"1003", x"0E73", x"0D19", x"0B3A", x"092A", x"078C", x"05AE", x"0398", x"021F", x"0091", x"FECD", x"FDFC", x"FDCD", x"FD82", x"FDBA", x"FE6D", x"FE6C", x"FEA8", x"FFEB", x"010B", x"01E1", x"034D", x"0405", x"03B7", x"0445", x"0545", x"054F", x"0555", x"056F", x"042D", x"02B7", x"02D4", x"0278", x"0070", x"FE44", x"FB7E", x"F802", x"F67A", x"F7A7", x"F927", x"FAD4", x"FD51", x"FF18", x"0026", x"01ED", x"035F", x"0377", x"036E", x"034F", x"026D", x"0210", x"025C", x"01D3", x"00B2", x"FF62", x"FCCB", x"F9B0", x"F7D4", x"F692", x"F57D", x"F5BB", x"F694", x"F720", x"F8D8", x"FBDB", x"FE64", x"00B9", x"030B", x"03E0", x"03C8", x"04A3", x"059D", x"061E", x"0768", x"08AE", x"08C3", x"0936", x"0A35", x"09C6", x"0811", x"062F", x"037F", x"0102", x"00FA", x"02C3", x"04CD", x"0750", x"098F", x"0A56", x"0AA8", x"0B1A", x"0B21", x"0B30", x"0BD6", x"0BFD", x"0BCE", x"0BFD", x"0BD3", x"0B2F", x"0AF5", x"0A58", x"08BF", x"07B0", x"078C", x"077F", x"0826", x"09A8", x"0A4C", x"0A54", x"0B14", x"0BAB", x"0B96", x"0BBF", x"0B32", x"08F7", x"0694", x"04BE", x"027C", x"00A9", x"FFBB", x"FE61", x"FCA0", x"FC0A", x"FB9F", x"FA4D", x"F8E6", x"F75B", x"F523", x"F42E", x"F5CE", x"F8D8", x"FC99", x"00FB", x"0480", x"068F", x"083B", x"098C", x"0A1D", x"0AC8", x"0B8A", x"0BA7", x"0B82", x"0B66", x"0A95", x"0926", x"07C4", x"05AF", x"0303", x"00E6", x"FF5E", x"FDF8", x"FD63", x"FDB4", x"FE05", x"FEBC", x"003F", x"018F", x"022D", x"02A0", x"0256", x"0143", x"00A8", x"00D1", x"013E", x"027B", x"047C", x"060F", x"0758", x"08E8", x"09BC", x"0931", x"083D", x"06CF", x"04F1", x"0442", x"0570", x"071D", x"08DD", x"0ACF", x"0C00", x"0C46", x"0C86", x"0C99", x"0BC2", x"0AA3", x"0967", x"079B", x"05A8", x"040F", x"0211", x"FFF5", x"FE31", x"FC5E", x"FAA4", x"F9F3", x"F9DB", x"F9E5", x"FA78", x"FB2B", x"FB70", x"FBFB", x"FD4A", x"FE82", x"FFD7", x"0182", x"0274", x"02D3", x"0392", x"0447", x"047F", x"0516", x"0597", x"0504", x"04A7", x"04F5", x"0450", x"029D", x"00A0", x"FD61", x"F9AF", x"F82E", x"F8F7", x"FA99", x"FD72", x"0102", x"0384", x"0592", x"0806", x"09A9", x"0A1D", x"0A7D", x"0A39", x"0938", x"08B1", x"086A", x"0765", x"0636", x"04C3", x"021B", x"FF4E", x"FD5B", x"FB7C", x"FA10", x"F9C5", x"F984", x"F8F2", x"F967", x"FA47", x"FA93", x"FB17", x"FB5D", x"FA2D", x"F8A1", x"F7D2", x"F687", x"F51A", x"F468", x"F2EC", x"F076", x"EEF4", x"EE0C", x"EC4F", x"EA94", x"E8E6", x"E60B", x"E3C9", x"E462", x"E6D6", x"EA50", x"EF32", x"F3E0", x"F70B", x"F9BC", x"FC4D", x"FDC8", x"FEF9", x"0068", x"014C", x"01C1", x"022B", x"01D5", x"00A6", x"FF83", x"FE11", x"FC57", x"FB8C", x"FB93", x"FBF3", x"FD4F", x"FF1B", x"0031", x"00FB", x"020A", x"02AC", x"0326", x"0429", x"0481", x"03D4", x"0322", x"0228", x"0071", x"FF1D", x"FE10", x"FC1D", x"FA1C", x"F8EE", x"F791", x"F5BF", x"F447", x"F25F", x"EFD2", x"EEDB", x"F044", x"F312", x"F72F", x"FC36", x"005A", x"0347", x"05BC", x"0763", x"07DE", x"082A", x"0843", x"07F8", x"07C1", x"07A7", x"06C8", x"056C", x"039B", x"00D6", x"FD86", x"FAAF", x"F819", x"F5F1", x"F4FB", x"F4A1", x"F443", x"F488", x"F582", x"F64B", x"F738", x"F87D", x"F905", x"F905", x"F981", x"FA19", x"FA86", x"FBCF", x"FD6F", x"FE6E", x"FFCE", x"01F8", x"035D", x"03CE", x"03D1", x"0279", x"0010", x"FF50", x"008C", x"0264", x"04F1", x"07E5", x"0963", x"09C8", x"0A66", x"0A6D", x"093D", x"080B", x"06E2", x"052C", x"03E8", x"031B", x"01BA", x"FFD8", x"FE09", x"FBB9", x"F94C", x"F79C", x"F62E", x"F4C0", x"F408", x"F385", x"F2EE", x"F320", x"F424", x"F528", x"F6A8", x"F872", x"F96B", x"FA1C", x"FB3B", x"FBEF", x"FC52", x"FD24", x"FD0E", x"FBB5", x"FADF", x"FA67", x"F91D", x"F7A8", x"F5AE", x"F174", x"EC8E", x"E9BD", x"E8A1", x"E908", x"EBDA", x"EF78", x"F20E", x"F4D7", x"F7E1", x"F9D2", x"FB1C", x"FC9E", x"FD5B", x"FDAE", x"FECB", x"FF8E", x"FFA5", x"FF95", x"FEB0", x"FC53", x"F9F9", x"F7D9", x"F574", x"F428", x"F406", x"F399", x"F386", x"F4BF", x"F60A", x"F784", x"FA27", x"FC3F", x"FCD0", x"FD8B", x"FE41", x"FDE8", x"FE1A", x"FEE8", x"FE1E", x"FCDC", x"FCD5", x"FCAE", x"FBD1", x"FB7C", x"F9E6", x"F5E3", x"F261", x"F100", x"F09A", x"F1F4", x"F52A", x"F7AD", x"F8DE", x"FA38", x"FB09", x"FAA0", x"FA63", x"FA4E", x"F9B5", x"F983", x"F9BF", x"F95B", x"F88A", x"F799", x"F5AF", x"F360", x"F1A9", x"F03E", x"EF82", x"F068", x"F1F2", x"F31D", x"F48F", x"F5AA", x"F5DF", x"F652", x"F742", x"F795", x"F7AA", x"F80C", x"F76F", x"F62C", x"F540", x"F3D1", x"F14F", x"EF60", x"EDF4", x"EC2A", x"EAC9", x"E9D7", x"E797", x"E4DE", x"E3DA", x"E49E", x"E732", x"EC27", x"F1DB", x"F644", x"F998", x"FC1D", x"FD43", x"FDE9", x"FEDE", x"FFB6", x"0092", x"01F3", x"0305", x"0356", x"0363", x"02B5", x"010F", x"FF7D", x"FE65", x"FD69", x"FD4C", x"FE20", x"FEB6", x"FEFA", x"FF7B", x"FFC2", x"FFAA", x"003E", x"00D1", x"00B9", x"00AD", x"00EA", x"00C2", x"010B", x"025C", x"034F", x"0403", x"057D", x"0740", x"0871", x"09CA", x"0A58", x"0871", x"0566", x"036E", x"0277", x"02D5", x"0518", x"0782", x"0831", x"0800", x"0779", x"058D", x"0302", x"00BE", x"FE57", x"FBEC", x"FA95", x"F9C0", x"F88C", x"F74F", x"F604", x"F463", x"F300", x"F26B", x"F224", x"F258", x"F32D", x"F433", x"F55E", x"F70A", x"F8DE", x"FAEA", x"FD88", x"0000", x"0200", x"03C1", x"04DD", x"051D", x"05AD", x"066D", x"063F", x"05D0", x"05C1", x"051E", x"042D", x"03CE", x"0239", x"FE5B", x"FA74", x"F7D0", x"F64E", x"F741", x"FAB4", x"FDEA", x"FFF7", x"01F1", x"0342", x"035E", x"03A9", x"0405", x"039E", x"034B", x"036F", x"0330", x"02A8", x"025B", x"0138", x"FF71", x"FD9D", x"FB60", x"F928", x"F819", x"F7B6", x"F73E", x"F759", x"F761", x"F6AF", x"F685", x"F73E", x"F781", x"F7A9", x"F842", x"F7C2", x"F675", x"F5DF", x"F4E3", x"F2A6", x"F0FF", x"F067", x"EF85", x"EF71", x"F02A", x"EEED", x"EB9E", x"E8E8", x"E746", x"E6E4", x"E958", x"EDD3", x"F1B5", x"F507", x"F84A", x"FA49", x"FB1D", x"FBBC", x"FC19", x"FC1F", x"FC9A", x"FD48", x"FD80", x"FD95", x"FD5A", x"FCD1", x"FC8E", x"FC83", x"FC8A", x"FD55", x"FF05", x"00C7", x"02A2", x"0498", x"0599", x"0613", x"0718", x"0837", x"091A", x"0A68", x"0B50", x"0ACE", x"09BF", x"0889", x"0622", x"0342", x"011B", x"FF15", x"FD33", x"FC74", x"FBCB", x"F9D8", x"F7B8", x"F695", x"F692", x"F89A", x"FD21", x"0256", x"06C0", x"0A3A", x"0C3E", x"0C82", x"0C0C", x"0B6B", x"0AB3", x"0A68", x"0A72", x"0A11", x"0905", x"075E", x"0491", x"00E8", x"FD57", x"FA0D", x"F736", x"F5C2", x"F52D", x"F48D", x"F3E8", x"F37E", x"F2EC", x"F2B4", x"F37D", x"F4C6", x"F61D", x"F7E4", x"F9B5", x"FB0D", x"FC74", x"FE08", x"FF29", x"0065", x"0278", x"04DD", x"074D", x"09F9", x"0B6C", x"0AB3", x"0901", x"07C3", x"0750", x"089D", x"0BD9", x"0EF9", x"10B2", x"1164", x"10E4", x"0EE3", x"0C83", x"0A3E", x"078A", x"04E3", x"02F9", x"012F", x"FF4C", x"FDCC", x"FC37", x"FA29", x"F869", x"F702", x"F588", x"F46B", x"F3F1", x"F3A1", x"F3CD", x"F4EF", x"F697", x"F8A8", x"FB49", x"FE27", x"00E0", x"038F", x"057B", x"0687", x"0728", x"0733", x"0680", x"05F8", x"0574", x"046F", x"0391", x"02F8", x"00C4", x"FCED", x"F92D", x"F5CD", x"F3C5", x"F513", x"F8EA", x"FC8D", x"FFA3", x"0250", x"0353", x"0353", x"0408", x"048B", x"045C", x"04CC", x"05C4", x"061B", x"0693", x"0717", x"063A", x"0456", x"0264", x"FFFE", x"FD5E", x"FBDA", x"FAFA", x"FA5E", x"FAC2", x"FBEC", x"FD22", x"FEE8", x"0134", x"033C", x"0546", x"0768", x"0892", x"0950", x"0A37", x"0A89", x"0A55", x"0AE1", x"0B8C", x"0BE4", x"0D25", x"0E6E", x"0D75", x"0AEA", x"084D", x"0575", x"03D2", x"055F", x"086F", x"0B01", x"0DA0", x"0FFE", x"10B3", x"10A4", x"109B", x"0FA7", x"0E28", x"0D94", x"0D58", x"0CD2", x"0C36", x"0B28", x"08F3", x"0677", x"0429", x"01E9", x"0020", x"FF1A", x"FE46", x"FDCC", x"FDAF", x"FD76", x"FD50", x"FDC0", x"FE58", x"FF46", x"00C9", x"01C7", x"019E", x"0103", x"FFB9", x"FD20", x"FA90", x"F89D", x"F672", x"F4DD", x"F4F0", x"F4C6", x"F321", x"F16A", x"F00B", x"EF11", x"F0DF", x"F5E6", x"FB79", x"0027", x"0458", x"06C6", x"0763", x"0813", x"0908", x"0950", x"09E4", x"0B37", x"0C0E", x"0C67", x"0CC2", x"0BFB", x"0A08", x"082C", x"0689", x"04F6", x"0460", x"0470", x"0410", x"038F", x"0352", x"02CD", x"0280", x"030F", x"03CE", x"04BA", x"0665", x"081B", x"0992", x"0B7E", x"0D5D", x"0E98", x"1025", x"1235", x"1402", x"1632", x"18FD", x"19F2", x"1873", x"15DB", x"12A3", x"0FB3", x"0FA1", x"1229", x"14A5", x"167D", x"17C6", x"1741", x"1580", x"143C", x"12EE", x"10FC", x"0F8F", x"0E9B", x"0D2B", x"0BDC", x"0AE7", x"094A", x"0768", x"05F8", x"0485", x"0308", x"022D", x"0174", x"00A1", x"0069", x"00B8", x"0142", x"02BC", x"04D6", x"0709", x"09AE", x"0C37", x"0D99", x"0E70", x"0F54", x"0F58", x"0EF9", x"0F13", x"0E3E", x"0C5A", x"0B55", x"0A83", x"0804", x"04DF", x"01D1", x"FE09", x"FBC1", x"FD63", x"00D7", x"0405", x"0766", x"09D9", x"0A16", x"0A4A", x"0B8C", x"0C36", x"0CB3", x"0E47", x"0FC6", x"10C4", x"1272", x"13C5", x"1352", x"1213", x"103D", x"0D39", x"0A04", x"0772", x"04B0", x"020A", x"001C", x"FE4E", x"FC82", x"FB66", x"FA80", x"F99A", x"F95B", x"F91E", x"F83C", x"F79B", x"F718", x"F5D0", x"F4B8", x"F42B", x"F308", x"F224", x"F2D6", x"F35D", x"F27D", x"F128", x"EF54", x"ECFC", x"ECE7", x"F058", x"F547", x"FAA5", x"0081", x"0529", x"07E4", x"0A2E", x"0BE3", x"0C45", x"0C42", x"0C8D", x"0C76", x"0C3E", x"0C42", x"0BE5", x"0B14", x"0A52", x"0959", x"0819", x"06FC", x"05C8", x"04A6", x"040E", x"03C4", x"0352", x"0372", x"03DA", x"0430", x"053D", x"06D5", x"076E", x"073C", x"06DA", x"052E", x"0237", x"FF94", x"FCB6", x"F914", x"F6F3", x"F6D2", x"F676", x"F59B", x"F4F8", x"F343", x"F177", x"F2E3", x"F754", x"FC60", x"01B9", x"066C", x"085E", x"085C", x"089A", x"0880", x"07E8", x"0848", x"093F", x"09B7", x"0A4A", x"0AF8", x"0A39", x"087B", x"068D", x"0425", x"0188", x"FFBA", x"FE29", x"FC60", x"FB15", x"FA12", x"F939", x"F91B", x"F9DF", x"FAE9", x"FC9C", x"FEBD", x"005E", x"01B6", x"0330", x"0408", x"04B6", x"0627", x"07BB", x"094B", x"0C13", x"0F67", x"1159", x"120D", x"11C1", x"0FD0", x"0E1B", x"0F0B", x"11D2", x"14DE", x"181B", x"1A48", x"1A27", x"1906", x"17F7", x"1642", x"1428", x"128F", x"10CC", x"0EA5", x"0CD0", x"0B0B", x"0915", x"0771", x"0641", x"04FE", x"03E1", x"02C2", x"0163", x"004C", x"FFB8", x"FF31", x"FF43", x"0017", x"010B", x"02AC", x"0543", x"0743", x"0810", x"088C", x"0827", x"0670", x"050A", x"03E8", x"0133", x"FE17", x"FC35", x"F9E3", x"F69E", x"F3AF", x"F009", x"EB14", x"E84A", x"E941", x"EBE9", x"EF9A", x"F444", x"F74D", x"F84E", x"F9A8", x"FB7C", x"FC8F", x"FE08", x"0063", x"022E", x"03C7", x"05C6", x"0709", x"06F0", x"0667", x"053F", x"030D", x"0087", x"FDE1", x"FB1A", x"F8F8", x"F7F9", x"F7C8", x"F87A", x"F9A1", x"FA98", x"FBA5", x"FCE4", x"FD8E", x"FDF0", x"FEAA", x"FEF7", x"FEB7", x"FEDB", x"FEAC", x"FD6F", x"FCAF", x"FD10", x"FD0F", x"FC5B", x"FB51", x"F8E6", x"F59A", x"F455", x"F5C7", x"F881", x"FC45", x"0078", x"0355", x"0493", x"054E", x"053A", x"0414", x"02D6", x"0219", x"0158", x"005A", x"FF27", x"FD72", x"FB61", x"F951", x"F77D", x"F5DE", x"F41E", x"F255", x"F156", x"F138", x"F16E", x"F22A", x"F36D", x"F44D", x"F52A", x"F717", x"F928", x"FA35", x"FB07", x"FB83", x"FA48", x"F83D", x"F661", x"F35D", x"EF74", x"ED2A", x"EC5F", x"EB57", x"EA80", x"E9C4", x"E755", x"E527", x"E628", x"E9DD", x"EE8E", x"F464", x"F9C0", x"FC91", x"FDEA", x"FF4C", x"FFBD", x"FFB8", x"00AC", x"0218", x"0365", x"0539", x"0728", x"080B", x"0853", x"0851", x"0791", x"067E", x"05B1", x"04AF", x"03A5", x"0318", x"027E", x"01ED", x"0213", x"028B", x"031D", x"0466", x"0604", x"06FE", x"0829", x"0985", x"0A14", x"0A37", x"0AC4", x"0ACD", x"0AB0", x"0BE0", x"0D65", x"0D6B", x"0C40", x"09C4", x"0582", x"01D3", x"00E5", x"01E7", x"03D1", x"0667", x"081A", x"07A9", x"065A", x"04CA", x"02C0", x"010B", x"004E", x"FFDB", x"FF7D", x"FF3F", x"FED1", x"FE33", x"FE15", x"FE1C", x"FE4E", x"FEAE", x"FEB7", x"FE61", x"FE7A", x"FED2", x"FF17", x"003F", x"0235", x"041C", x"06CE", x"0A47", x"0CDA", x"0E7C", x"1030", x"10DB", x"1045", x"0FDE", x"0ED5", x"0BD7", x"08D0", x"06CD", x"045C", x"01BC", x"FFA6", x"FC2A", x"F75C", x"F475", x"F410", x"F4E2", x"F76A", x"FABB", x"FC1B", x"FC01", x"FC57", x"FC89", x"FC89", x"FDBB", x"FF5F", x"004A", x"0181", x"0305", x"0395", x"0380", x"0358", x"0209", x"FFD8", x"FD84", x"FA92", x"F6E9", x"F3B6", x"F0ED", x"EE63", x"ECF4", x"EC53", x"EBAA", x"EB59", x"EB6D", x"EB01", x"EAB2", x"EB22", x"EB54", x"EB27", x"EB27", x"EA6E", x"E8AA", x"E7A1", x"E795", x"E753", x"E728", x"E6E3", x"E53D", x"E35A", x"E3A1", x"E645", x"EA6E", x"F04E", x"F65A", x"FABE", x"FDCD", x"0049", x"018B", x"01F9", x"0263", x"0292", x"025F", x"0254", x"0256", x"0221", x"0220", x"0249", x"025F", x"026F", x"024D", x"01D0", x"01DC", x"026C", x"0317", x"0400", x"0525", x"05AC", x"061D", x"078C", x"08E8", x"09E5", x"0B4C", x"0C7F", x"0C3C", x"0BA1", x"0ABC", x"07FB", x"0482", x"027B", x"012C", x"FFF9", x"FFE4", x"FF49", x"FC92", x"FA24", x"FA1B", x"FB86", x"FE68", x"02BE", x"059C", x"058E", x"0482", x"02F8", x"0074", x"FE9B", x"FE02", x"FD48", x"FCB8", x"FD2D", x"FD5C", x"FCC9", x"FC49", x"FB35", x"F91C", x"F72D", x"F588", x"F389", x"F20F", x"F132", x"F005", x"EF3A", x"EF73", x"EFE8", x"F0C2", x"F2B0", x"F479", x"F5BC", x"F79C", x"F9A3", x"FAEC", x"FCAB", x"FEA2", x"FF9B", x"00C2", x"0344", x"05A5", x"0746", x"08AF", x"0820", x"055F", x"0331", x"02EA", x"03CE", x"0642", x"098D", x"0AE3", x"09F7", x"0818", x"0518", x"0166", x"FE94", x"FC59", x"FA0C", x"F83F", x"F6CC", x"F4FD", x"F3AB", x"F303", x"F257", x"F1E2", x"F1C1", x"F0EF", x"EFF7", x"EFA2", x"EF2A", x"EEBA", x"EF74", x"F0B7", x"F215", x"F4F7", x"F88F", x"FB1A", x"FD5C", x"FF82", x"0000", x"FFCE", x"0043", x"FF83", x"FD17", x"FB25", x"F952", x"F699", x"F4B2", x"F31B", x"EF6C", x"EAF8", x"E86E", x"E75A", x"E817", x"EB9A", x"EF77", x"F127", x"F219", x"F2E4", x"F302", x"F3DC", x"F633", x"F830", x"F9A3", x"FB61", x"FC9B", x"FD21", x"FE11", x"FED0", x"FE6B", x"FD9B", x"FC32", x"F990", x"F6F5", x"F4F9", x"F31A", x"F1FC", x"F23C", x"F2D0", x"F3B5", x"F5BC", x"F7C7", x"F937", x"FB0C", x"FCC1", x"FD6E", x"FE28", x"FF01", x"FE7B", x"FD68", x"FD2C", x"FD20", x"FD3B", x"FE57", x"FEF0", x"FDC9", x"FC7C", x"FC66", x"FD54", x"FFF4", x"0436", x"07CC", x"09A9", x"0A6B", x"09E3", x"084B", x"06B7", x"0558", x"03B5", x"0208", x"002F", x"FDD7", x"FB71", x"F965", x"F768", x"F5AD", x"F441", x"F272", x"F0C4", x"F00F", x"EFF5", x"F043", x"F170", x"F29A", x"F325", x"F444", x"F644", x"F83E", x"FA81", x"FD54", x"FF29", x"FFDC", x"0082", x"003D", x"FE38", x"FC0D", x"FA70", x"F8CA", x"F7F8", x"F880", x"F840", x"F6CE", x"F5FD", x"F657", x"F7B2", x"FB16", x"FFB0", x"02E6", x"044F", x"04B0", x"03C9", x"023C", x"01A7", x"01CC", x"01FB", x"0298", x"036C", x"037B", x"033E", x"02F4", x"0218", x"00FB", x"0035", x"FF71", x"FEAF", x"FE93", x"FE67", x"FDD0", x"FD38", x"FC89", x"FB6B", x"FADC", x"FB27", x"FB96", x"FCAF", x"FEA3", x"006F", x"01FE", x"03F6", x"0561", x"05CC", x"0688", x"0771", x"079E", x"07A3", x"0731", x"04B2", x"00E2", x"FE08", x"FC76", x"FC98", x"FF46", x"02B6", x"0494", x"04E2", x"0413", x"01BC", x"FF3D", x"FDD5", x"FCE1", x"FC3B", x"FC5B", x"FCA8", x"FC94", x"FCE2", x"FD60", x"FD97", x"FE0A", x"FE84", x"FE6A", x"FE2B", x"FE1B", x"FDCD", x"FDCA", x"FE8F", x"FF5F", x"007E", x"02AF", x"051F", x"0781", x"0A5D", x"0CDB", x"0DE2", x"0EB3", x"0F37", x"0E31", x"0C63", x"0AEA", x"08B2", x"0628", x"04B9", x"02FC", x"FF73", x"FBE4", x"F969", x"F7BD", x"F87A", x"FBFF", x"FF87", x"019C", x"0330", x"03FA", x"040E", x"051F", x"073C", x"08FC", x"0A86", x"0C2D", x"0CFC", x"0D35", x"0D51", x"0CEE", x"0BCF", x"0A54", x"080D", x"04CB", x"0136", x"FD48", x"F946", x"F5E0", x"F2DA", x"EFD7", x"EDBD", x"ECB5", x"EC30", x"ECA0", x"EE15", x"EF06", x"EF68", x"F040", x"F093", x"EFC5", x"EF0C", x"EE93", x"EDA3", x"ED7A", x"EECD", x"EF82", x"EF3B", x"EF69", x"F086", x"F2B0", x"F75C", x"FDEB", x"03EC", x"0889", x"0C42", x"0E82", x"0F4D", x"0F96", x"0F6B", x"0E71", x"0D1F", x"0BED", x"0A95", x"0915", x"07C5", x"06F4", x"067B", x"061A", x"057E", x"04A5", x"038D", x"023F", x"0177", x"00F4", x"0021", x"FF16", x"FECC", x"FF11", x"0018", x"025A", x"050D", x"06A4", x"0763", x"0792", x"0636", x"0360", x"009A", x"FDED", x"FB70", x"FA7B", x"FAFF", x"FB02", x"FA5F", x"FA68", x"FB2B", x"FCB4", x"FFF8", x"03E9", x"0647", x"06F9", x"06E7", x"05C1", x"040D", x"033B", x"035A", x"03EB", x"0542", x"0715", x"0848", x"088B", x"0840", x"0762", x"0634", x"0503", x"03CD", x"02B6", x"01EA", x"0151", x"00FC", x"00D5", x"0051", x"FF8F", x"FF57", x"FF82", x"FFFC", x"017A", x"03A3", x"056A", x"0763", x"09AB", x"0AE7", x"0B30", x"0BEC", x"0CBE", x"0D74", x"0F36", x"111D", x"10FC", x"0FC1", x"0F26", x"0F02", x"100F", x"1342", x"1671", x"177C", x"1715", x"15AF", x"12C1", x"0FBE", x"0DC8", x"0C0E", x"0A9B", x"0A20", x"09DD", x"0923", x"087A", x"07AB", x"0663", x"0535", x"041A", x"02A5", x"0143", x"0008", x"FE8A", x"FD54", x"FC9C", x"FBD7", x"FB92", x"FC64", x"FD89", x"FEE2", x"00F8", x"0299", x"0331", x"03DB", x"042E", x"030A", x"017F", x"003E", x"FE51", x"FC99", x"FC23", x"FB13", x"F844", x"F57A", x"F340", x"F1B6", x"F2CD", x"F68E", x"FA56", x"FD28", x"FFB7", x"013C", x"020B", x"03BE", x"061C", x"0839", x"0A8B", x"0CEF", x"0EA6", x"0FF5", x"1115", x"117C", x"113B", x"1065", x"0E64", x"0BB3", x"08FF", x"064C", x"03FE", x"02C4", x"01B1", x"007F", x"0034", x"0096", x"0102", x"023D", x"03EE", x"0470", x"0489", x"0539", x"054A", x"0466", x"03E2", x"0308", x"014C", x"00A8", x"0145", x"00F1", x"FFC7", x"FF20", x"FEA5", x"FF0D", x"023E", x"0712", x"0B03", x"0DF1", x"0FE4", x"1009", x"0F03", x"0E00", x"0C93", x"0A70", x"0849", x"0613", x"0369", x"009D", x"FE07", x"FBE9", x"FA76", x"F9AB", x"F923", x"F8E6", x"F8BD", x"F89E", x"F8EB", x"F972", x"F953", x"F8F2", x"F902", x"F959", x"FA66", x"FCE2", x"FFBF", x"01D7", x"03A9", x"04EC", x"0469", x"029D", x"0088", x"FDDD", x"FB21", x"FA18", x"FA12", x"F96D", x"F88B", x"F81C", x"F7CC", x"F88C", x"FB6B", x"FF1F", x"01ED", x"0424", x"05A2", x"05E4", x"059D", x"05A7", x"05C9", x"0607", x"06BE", x"07A1", x"0810", x"082B", x"0831", x"0877", x"0932", x"0A2C", x"0B26", x"0C39", x"0CFF", x"0D6A", x"0DBB", x"0D7B", x"0C08", x"0A15", x"0862", x"06B5", x"05AC", x"0622", x"0722", x"0835", x"0A29", x"0C57", x"0D37", x"0D5D", x"0D43", x"0BFA", x"0A5E", x"09C9", x"08CF", x"0643", x"0391", x"0187", x"0005", x"00DF", x"0475", x"0819", x"0A32", x"0B34", x"0A55", x"07B7", x"0532", x"0371", x"01CD", x"00FB", x"016A", x"0217", x"02EB", x"041B", x"050C", x"058F", x"0634", x"06B1", x"06F6", x"0783", x"083E", x"08A9", x"0943", x"09BC", x"09A9", x"09C7", x"0A83", x"0B64", x"0D0B", x"0FA2", x"11FE", x"13DF", x"15B2", x"162E", x"14C9", x"1283", x"0F5B", x"0AFB", x"0745", x"04E1", x"021D", x"FF03", x"FC6F", x"F9D1", x"F7C6", x"F85D", x"FADD", x"FD21", x"FF04", x"005D", x"0048", x"FFF1", x"00D0", x"0256", x"0429", x"06B9", x"0946", x"0B21", x"0CB5", x"0DE3", x"0E34", x"0E0A", x"0D45", x"0B44", x"0897", x"0580", x"01FC", x"FEC8", x"FC47", x"F9C6", x"F789", x"F654", x"F5AE", x"F5A0", x"F6F7", x"F875", x"F8E5", x"F91C", x"F923", x"F7E1", x"F642", x"F509", x"F2F5", x"F071", x"EFBD", x"F00F", x"F003", x"F046", x"F0E0", x"F0D4", x"F206", x"F63F", x"FBEE", x"015E", x"068E", x"0A5F", x"0BC7", x"0C15", x"0C1B", x"0B45", x"09EA", x"0909", x"0848", x"076D", x"06C4", x"0650", x"05DF", x"05AF", x"05B4", x"05A7", x"0560", x"04BE", x"0411", x"03CB", x"03A5", x"0354", x"0320", x"02ED", x"02AF", x"035F", x"054D", x"075A", x"0927", x"0AD1", x"0B47", x"09F8", x"07EE", x"0529", x"015D", x"FE08", x"FC88", x"FBF4", x"FBAD", x"FC16", x"FC90", x"FC9F", x"FDB5", x"0032", x"028F", x"03EC", x"0491", x"0408", x"0254", x"00BB", x"FFC8", x"FF2C", x"FF1D", x"FFD9", x"009F", x"00C8", x"004B", x"FF4D", x"FE1C", x"FD2B", x"FCA0", x"FC70", x"FC5B", x"FC4A", x"FC53", x"FCA2", x"FCCC", x"FC8E", x"FC31", x"FBCA", x"FB60", x"FBE3", x"FD8B", x"FFA6", x"020C", x"04CD", x"06CD", x"0783", x"07B2", x"0756", x"0644", x"05F7", x"0717", x"082B", x"088B", x"08BF", x"0824", x"0705", x"0761", x"0950", x"0B05", x"0BFF", x"0C76", x"0B3E", x"08DA", x"06CA", x"04FC", x"02D4", x"013E", x"0061", x"FF57", x"FE7F", x"FE17", x"FD54", x"FC45", x"FB89", x"FAE8", x"FA39", x"FA21", x"FA4E", x"FA44", x"FA67", x"FA8C", x"FA6D", x"FA2A", x"FA0B", x"F9E2", x"FA34", x"FB82", x"FD6B", x"0002", x"02F0", x"0521", x"064E", x"06A4", x"058F", x"0341", x"0117", x"FF09", x"FC3A", x"F94D", x"F651", x"F29D", x"EFAF", x"EF75", x"F107", x"F351", x"F65B", x"F8D7", x"F9B6", x"FA5C", x"FBC8", x"FCFB", x"FE4C", x"0054", x"020F", x"032A", x"0484", x"0581", x"055D", x"04C3", x"03E0", x"0244", x"0095", x"FF53", x"FDF6", x"FC9E", x"FBA5", x"FAB5", x"F9A2", x"F8D4", x"F811", x"F7DD", x"F8B3", x"FA72", x"FCA3", x"FF61", x"01C7", x"0310", x"03FA", x"0448", x"0310", x"018F", x"0105", x"00B3", x"0084", x"0133", x"0187", x"00CD", x"0142", x"0401", x"0781", x"0B57", x"0F3B", x"111B", x"107A", x"0F2C", x"0D59", x"0A4F", x"06EE", x"03F4", x"0093", x"FD38", x"FA92", x"F83F", x"F5CF", x"F41F", x"F33C", x"F2B7", x"F25C", x"F22D", x"F1D0", x"F155", x"F101", x"F0FC", x"F0FA", x"F0CA", x"F0BA", x"F189", x"F350", x"F5D2", x"F925", x"FC78", x"FEA0", x"FF98", x"FFEE", x"FEE4", x"FC78", x"FA5F", x"F8F3", x"F7A7", x"F6FC", x"F6F3", x"F626", x"F4D7", x"F4F4", x"F699", x"F874", x"FA94", x"FC4F", x"FC4D", x"FAE7", x"F9A3", x"F839", x"F655", x"F4DD", x"F41B", x"F360", x"F2EB", x"F2F3", x"F2E3", x"F2A6", x"F30D", x"F409", x"F534", x"F69B", x"F809", x"F907", x"F9C0", x"FA4F", x"FA8E", x"FA52", x"F9D3", x"F91E", x"F8EB", x"F99D", x"FB64", x"FE3D", x"01A0", x"047C", x"064C", x"0710", x"063F", x"0424", x"022B", x"00E3", x"FFA8", x"FEFE", x"FED4", x"FE25", x"FD93", x"FEC4", x"0126", x"033C", x"0503", x"05D3", x"046A", x"0209", x"002F", x"FE59", x"FC94", x"FC25", x"FCA9", x"FD83", x"FF5A", x"01D9", x"03B3", x"050C", x"0664", x"0700", x"073D", x"07CB", x"082B", x"07EF", x"07B6", x"075C", x"0684", x"05AF", x"050E", x"0458", x"0437", x"0533", x"071F", x"09D3", x"0CA0", x"0E57", x"0EA2", x"0D83", x"0A97", x"06D9", x"03CB", x"016F", x"FFAA", x"FF11", x"FE73", x"FC97", x"FB24", x"FB42", x"FC17", x"FD9A", x"0004", x"013E", x"00BF", x"0086", x"00C4", x"00B9", x"016B", x"02FA", x"03E5", x"0480", x"05C4", x"063B", x"0562", x"041D", x"01E0", x"FE63", x"FB07", x"F847", x"F54F", x"F298", x"F0AB", x"EED4", x"ED34", x"EC41", x"EB60", x"EA7F", x"EA2B", x"EA5E", x"EAF1", x"EBF1", x"EC6F", x"EC12", x"EB64", x"EA10", x"E7C5", x"E5FE", x"E54D", x"E519", x"E618", x"E86F", x"EA00", x"EABC", x"ECBB", x"F037", x"F472", x"FA08", x"FFC9", x"0322", x"0451", x"04E4", x"043F", x"0291", x"0156", x"0043", x"FEB2", x"FD8B", x"FCED", x"FBC0", x"FA1B", x"F8B9", x"F746", x"F5F5", x"F55F", x"F542", x"F521", x"F528", x"F559", x"F573", x"F55F", x"F4E7", x"F445", x"F403", x"F485", x"F60A", x"F8BA", x"FB90", x"FD60", x"FE6B", x"FE9C", x"FD06", x"FA3F", x"F7B2", x"F530", x"F31D", x"F299", x"F2FF", x"F285", x"F209", x"F2DE", x"F478", x"F6B7", x"F9F0", x"FCB0", x"FD86", x"FD96", x"FDCA", x"FD8E", x"FD2B", x"FD68", x"FD7A", x"FD0E", x"FCB1", x"FC59", x"FB50", x"FA30", x"F994", x"F94D", x"F98C", x"FAA4", x"FBF7", x"FD03", x"FDEB", x"FEA0", x"FED5", x"FEBB", x"FE55", x"FD9F", x"FCF5", x"FD01", x"FE0B", x"0027", x"02E2", x"0564", x"0742", x"083C", x"07E6", x"06E0", x"0655", x"065E", x"06E4", x"0832", x"0958", x"0925", x"08A7", x"092B", x"0A59", x"0C13", x"0E9D", x"107B", x"1098", x"1025", x"0F9C", x"0E45", x"0CD2", x"0C0E", x"0B46", x"0A80", x"0A8C", x"0AAA", x"09F0", x"08FA", x"07B7", x"059B", x"0396", x"0229", x"0093", x"FEE2", x"FD97", x"FC05", x"F9F7", x"F824", x"F624", x"F3B1", x"F1BD", x"F10E", x"F1BA", x"F43E", x"F809", x"FBC9", x"FEC8", x"0074", x"FFFC", x"FE32", x"FC02", x"F97E", x"F72B", x"F5CF", x"F3FE", x"F139", x"EF4A", x"EED5", x"EF77", x"F22F", x"F678", x"F9A1", x"FB6F", x"FD22", x"FE08", x"FE12", x"FEDF", x"FFCB", x"FFC4", x"FFF2", x"00B3", x"0078", x"FF8F", x"FEB4", x"FCA4", x"F9DC", x"F820", x"F720", x"F618", x"F5BE", x"F59E", x"F480", x"F33A", x"F256", x"F12A", x"F021", x"F049", x"F16F", x"F3C0", x"F745", x"FAB0", x"FD0D", x"FE66", x"FDF6", x"FBF7", x"F9EF", x"F852", x"F70F", x"F76C", x"F8E3", x"F949", x"F901", x"F983", x"FA68", x"FC28", x"FFD8", x"0388", x"04F3", x"04FD", x"0432", x"01DB", x"FF11", x"FD2C", x"FB10", x"F8F7", x"F802", x"F7AD", x"F6F2", x"F668", x"F5E9", x"F4B7", x"F39D", x"F312", x"F27A", x"F1BD", x"F143", x"F0AD", x"F008", x"EFCA", x"EFB0", x"EFA5", x"F010", x"F116", x"F2FD", x"F614", x"F967", x"FC0D", x"FE20", x"FF0E", x"FE21", x"FC5B", x"FA94", x"F879", x"F703", x"F76E", x"F82F", x"F80F", x"F822", x"F8DF", x"F9EF", x"FC5E", x"0037", x"031C", x"03EC", x"03B9", x"028B", x"007D", x"FEEF", x"FE7B", x"FE5F", x"FED4", x"0048", x"01C2", x"02CD", x"03E4", x"04E5", x"05B4", x"0705", x"08F4", x"0AF3", x"0CEB", x"0EBC", x"0FC9", x"0FF4", x"0F8B", x"0E5F", x"0C72", x"0A73", x"08DA", x"083E", x"090C", x"0AF5", x"0D0B", x"0EBA", x"0F2A", x"0DC8", x"0B46", x"089C", x"0639", x"04F6", x"0552", x"0601", x"0607", x"060D", x"068E", x"0714", x"0843", x"09F2", x"0A7D", x"0965", x"0801", x"066B", x"0476", x"0356", x"034C", x"03B1", x"04C7", x"0701", x"0936", x"0B09", x"0CCC", x"0E1D", x"0EA5", x"0F58", x"1030", x"109A", x"1121", x"119E", x"1184", x"1110", x"10D4", x"1027", x"0F01", x"0E35", x"0DE6", x"0E68", x"1054", x"12F2", x"1505", x"162D", x"15A0", x"1336", x"0FDD", x"0C95", x"0952", x"072F", x"0620", x"0490", x"023A", x"0079", x"FF41", x"FF0B", x"0132", x"0492", x"06EA", x"0859", x"0956", x"08E4", x"07E2", x"07C6", x"07A6", x"0735", x"07AE", x"0860", x"0828", x"07B2", x"06B5", x"041C", x"00DF", x"FE76", x"FC46", x"FAD2", x"FAEF", x"FB5F", x"FB52", x"FBA3", x"FBD3", x"FAD6", x"F959", x"F7D5", x"F5F6", x"F4DD", x"F53E", x"F602", x"F6AF", x"F710", x"F5FF", x"F392", x"F13B", x"EF12", x"ED8B", x"EDF7", x"EF55", x"EFE8", x"F04E", x"F16C", x"F2ED", x"F60E", x"FBB4", x"016D", x"0595", x"08C1", x"0AAD", x"0AD3", x"0AE0", x"0B72", x"0B92", x"0BB7", x"0C83", x"0CF4", x"0C9B", x"0C2B", x"0B48", x"09EA", x"0958", x"09B7", x"0A88", x"0BEB", x"0D90", x"0E72", x"0EC9", x"0ED8", x"0E43", x"0D48", x"0C6C", x"0BB9", x"0BA1", x"0CC7", x"0E61", x"0FF9", x"114A", x"1172", x"0FB8", x"0D27", x"0A14", x"0675", x"03DA", x"02E3", x"020A", x"00A8", x"FFBA", x"FF13", x"FF15", x"0175", x"05E1", x"09E0", x"0CC1", x"0E9F", x"0EAE", x"0D3B", x"0BCA", x"0A51", x"086C", x"06D0", x"05AD", x"043E", x"02CE", x"01C6", x"00CB", x"000F", x"002C", x"00CA", x"01A9", x"032C", x"04D5", x"061C", x"0729", x"081E", x"0853", x"081A", x"07BC", x"0737", x"0710", x"0827", x"0A38", x"0CCA", x"0F78", x"1148", x"1162", x"1067", x"0ED8", x"0CDE", x"0B9C", x"0B59", x"0AC2", x"095A", x"0826", x"0739", x"06CF", x"0827", x"0A96", x"0C10", x"0C46", x"0C0A", x"0AD4", x"0922", x"0869", x"088D", x"08EA", x"0A0D", x"0BC3", x"0CBA", x"0CCE", x"0C43", x"0AA9", x"0850", x"061F", x"03F1", x"01D1", x"0048", x"FF0A", x"FDA7", x"FC8B", x"FBAE", x"FA60", x"F912", x"F82D", x"F7B5", x"F8B0", x"FBBB", x"001F", x"04EE", x"0956", x"0BB4", x"0B92", x"09C9", x"06B8", x"02F5", x"0056", x"FE91", x"FC53", x"F9F2", x"F81D", x"F666", x"F616", x"F8B8", x"FC83", x"FFB7", x"029F", x"04A3", x"04D0", x"048E", x"04DC", x"04B9", x"04AE", x"05BB", x"06C6", x"073E", x"07B8", x"0777", x"05D0", x"040A", x"0260", x"006B", x"FF22", x"FED0", x"FE30", x"FD79", x"FD63", x"FD05", x"FC54", x"FC32", x"FC1A", x"FBE0", x"FCDB", x"FF2B", x"01B9", x"04C4", x"077C", x"0851", x"07C1", x"06C8", x"053A", x"0414", x"04C6", x"05B6", x"0575", x"04DC", x"03F2", x"02AA", x"031C", x"05EA", x"0894", x"0A0B", x"0AAB", x"0975", x"065D", x"0363", x"00D7", x"FE6B", x"FD21", x"FD4E", x"FDB6", x"FE03", x"FE21", x"FD44", x"FBA9", x"FA1E", x"F882", x"F714", x"F678", x"F64F", x"F627", x"F680", x"F6F5", x"F70A", x"F73A", x"F7AD", x"F7F4", x"F8D4", x"FAE4", x"FD75", x"0066", x"03A6", x"05CC", x"0640", x"05E8", x"049A", x"02A3", x"01BD", x"023C", x"0261", x"021A", x"01C6", x"00D6", x"0029", x"01CF", x"04CA", x"0720", x"087C", x"0881", x"065B", x"031C", x"0062", x"FDF6", x"FC0C", x"FB59", x"FB6A", x"FB6A", x"FBC9", x"FC68", x"FD04", x"FE45", x"0044", x"0262", x"04C4", x"077B", x"099F", x"0ADB", x"0BA7", x"0B88", x"0A5B", x"0900", x"0775", x"0586", x"042B", x"0412", x"04E3", x"0692", x"08E4", x"0A57", x"0A57", x"0999", x"07F8", x"0614", x"055A", x"0582", x"0516", x"03F9", x"0267", x"FFF9", x"FDCA", x"FD98", x"FE55", x"FEA0", x"FEC4", x"FE87", x"FD24", x"FBBA", x"FB46", x"FB42", x"FBB5", x"FD63", x"FF9A", x"0189", x"0378", x"0532", x"0666", x"0792", x"08D9", x"09D2", x"0AC9", x"0BDB", x"0CA3", x"0D24", x"0DC4", x"0DE8", x"0D6A", x"0CAC", x"0B52", x"0987", x"086D", x"0860", x"091A", x"0AE9", x"0CBC", x"0D5B", x"0CA1", x"0AE4", x"07C7", x"049F", x"02E9", x"01D4", x"008E", x"FFB4", x"FEC5", x"FD6F", x"FDDA", x"00C6", x"042F", x"072B", x"09A4", x"0A46", x"08AF", x"06BB", x"04B4", x"0206", x"FFCA", x"FE82", x"FD2A", x"FBCE", x"FAA3", x"F8E9", x"F69D", x"F4A1", x"F2BC", x"F114", x"F07F", x"F0C5", x"F140", x"F250", x"F382", x"F3C2", x"F354", x"F259", x"F040", x"EDE5", x"EC9A", x"EC38", x"ECD3", x"EEAE", x"F04E", x"F08C", x"EFFC", x"EEB2", x"ECC6", x"EC19", x"ED72", x"EF34", x"F0AF", x"F23E", x"F2CF", x"F31A", x"F551", x"F994", x"FDD3", x"01C6", x"04FF", x"0615", x"0579", x"0494", x"034B", x"0189", x"0050", x"FFA3", x"FEC1", x"FDB8", x"FC8A", x"FB1B", x"F9F7", x"F965", x"F92A", x"F95B", x"FA00", x"FA9C", x"FB63", x"FC8C", x"FD6A", x"FDD7", x"FE42", x"FE45", x"FDA8", x"FD51", x"FD5E", x"FD70", x"FDF1", x"FEA2", x"FE3D", x"FC9E", x"FA5C", x"F71D", x"F3BD", x"F1E1", x"F14F", x"F0CB", x"F053", x"EFC4", x"EE8A", x"EE4C", x"F0CF", x"F543", x"FA07", x"FEAA", x"01BA", x"0227", x"00DD", x"FEF5", x"FC95", x"FA54", x"F937", x"F8E5", x"F8DC", x"F932", x"F99C", x"F9FD", x"FAAF", x"FBA7", x"FC91", x"FD99", x"FECA", x"FFB2", x"00A6", x"01D2", x"02B3", x"0348", x"03D3", x"03E3", x"0346", x"02D7", x"0308", x"03E7", x"05C8", x"082A", x"09C4", x"0A43", x"09B5", x"0805", x"0605", x"0501", x"0480", x"03E0", x"0345", x"025D", x"00D3", x"0040", x"0199", x"03B5", x"05B5", x"078D", x"0858", x"07AB", x"06F6", x"06D5", x"06BF", x"06FA", x"07E0", x"084C", x"07AF", x"0661", x"0436", x"0162", x"FEBF", x"FC7B", x"FA30", x"F812", x"F5F6", x"F38E", x"F13A", x"EF5C", x"EDBB", x"EC4A", x"EB5D", x"EA5D", x"E988", x"E9A6", x"EAF2", x"ED49", x"F095", x"F3BD", x"F596", x"F617", x"F539", x"F312", x"F12A", x"F074", x"F034", x"F00F", x"F02B", x"EF86", x"EE70", x"EF30", x"F245", x"F63D", x"FAA5", x"FEF7", x"0143", x"0189", x"0159", x"006F", x"FE7A", x"FCB5", x"FB8F", x"FA42", x"F922", x"F881", x"F799", x"F670", x"F5A8", x"F4E7", x"F3F0", x"F325", x"F265", x"F1A8", x"F1A4", x"F263", x"F359", x"F496", x"F589", x"F595", x"F52D", x"F530", x"F5CD", x"F796", x"FAB0", x"FDCC", x"000E", x"016D", x"0150", x"FFE0", x"FEE4", x"FE99", x"FDFD", x"FD15", x"FBC7", x"F908", x"F61B", x"F54E", x"F642", x"F798", x"F955", x"FA7A", x"F99F", x"F7B3", x"F62F", x"F486", x"F2FE", x"F2C0", x"F35E", x"F402", x"F4AA", x"F507", x"F495", x"F3E8", x"F384", x"F336", x"F329", x"F358", x"F365", x"F36E", x"F3C5", x"F3BE", x"F360", x"F2ED", x"F210", x"F0A6", x"EFB2", x"EF6B", x"EFC0", x"F137", x"F38D", x"F554", x"F651", x"F69C", x"F5D5", x"F4CD", x"F52F", x"F67D", x"F7C8", x"F8F5", x"F94F", x"F81F", x"F738", x"F84B", x"FA94", x"FD5D", x"0075", x"0244", x"01CD", x"003D", x"FE37", x"FB77", x"F8DA", x"F74F", x"F650", x"F5D5", x"F64B", x"F756", x"F8F6", x"FB79", x"FE70", x"0114", x"0371", x"0500", x"0583", x"058F", x"0574", x"04D0", x"0407", x"0365", x"0238", x"004A", x"FE92", x"FD06", x"FC09", x"FC3E", x"FD52", x"FE22", x"FE9B", x"FE9F", x"FDD3", x"FD28", x"FD5B", x"FD78", x"FD27", x"FC4C", x"FA28", x"F6F6", x"F4F0", x"F4E4", x"F60B", x"F863", x"FB23", x"FC88", x"FC7B", x"FC65", x"FC1A", x"FBA7", x"FC00", x"FD0B", x"FDCD", x"FE93", x"FF73", x"FFD3", x"0026", x"0119", x"022A", x"0318", x"0435", x"04D3", x"04A4", x"046D", x"0463", x"0421", x"042C", x"044D", x"03B0", x"027F", x"017D", x"00F1", x"012A", x"0276", x"03D1", x"0475", x"044F", x"0310", x"0119", x"FFC6", x"FF7F", x"FFAF", x"008D", x"0164", x"00D6", x"FF9B", x"FF81", x"0067", x"01ED", x"044B", x"062D", x"05E0", x"0454", x"027C", x"FFDD", x"FCD0", x"FA6A", x"F83A", x"F5EF", x"F461", x"F394", x"F2DB", x"F2E0", x"F3C8", x"F4F5", x"F62C", x"F76A", x"F805", x"F819", x"F85F", x"F8CC", x"F95F", x"FA43", x"FAC5", x"FA5A", x"F964", x"F834", x"F713", x"F6CA", x"F752", x"F7C2", x"F7FB", x"F7BB", x"F674", x"F4F2", x"F4BE", x"F58F", x"F6E5", x"F8DA", x"FA11", x"F95B", x"F879", x"F93C", x"FB39", x"FE5E", x"02B0", x"064E", x"07F0", x"0904", x"09E5", x"09C3", x"0940", x"090D", x"0877", x"0782", x"06F0", x"066F", x"05CD", x"05B6", x"064D", x"06F8", x"07CE", x"0867", x"0878", x"087D", x"08D0", x"091B", x"0986", x"0A05", x"09BC", x"0898", x"073C", x"0581", x"03CE", x"02E8", x"0271", x"016B", x"FFF2", x"FDBD", x"FA66", x"F752", x"F5CE", x"F55C", x"F5AC", x"F6A4", x"F6C3", x"F594", x"F520", x"F671", x"F8FC", x"FCE5", x"016F", x"0463", x"0517", x"04A5", x"02F5", x"0024", x"FD8C", x"FB83", x"F99B", x"F85F", x"F806", x"F805", x"F8D9", x"FAA8", x"FC99", x"FE68", x"0008", x"00D4", x"00D2", x"0122", x"016E", x"016E", x"0201", x"0309", x"0375", x"039B", x"03FB", x"03EE", x"0423", x"0592", x"0766", x"08AB", x"097E", x"0943", x"079D", x"0620", x"0573", x"04E5", x"049F", x"043B", x"0250", x"FF47", x"FD40", x"FC80", x"FD22", x"FFCD", x"0330", x"056B", x"06E4", x"082E", x"0895", x"08A1", x"0910", x"08ED", x"07F5", x"06EA", x"058E", x"03A4", x"0240", x"017F", x"00A3", x"0031", x"0021", x"FF6E", x"FE44", x"FD69", x"FC5C", x"FB6D", x"FB83", x"FC3C", x"FCA9", x"FD35", x"FDE3", x"FE77", x"FFA8", x"01A6", x"0367", x"04A8", x"053E", x"04A1", x"0382", x"0312", x"0314", x"0379", x"048A", x"04CF", x"0320", x"00FD", x"FF9C", x"FF2C", x"00C6", x"0489", x"07DE", x"0996", x"0A80", x"0A6B", x"0906", x"07C7", x"06C6", x"04F5", x"0319", x"020E", x"0135", x"00BB", x"016E", x"0263", x"02DB", x"0362", x"036C", x"0260", x"0143", x"0097", x"001B", x"0046", x"0182", x"028D", x"030E", x"035B", x"0349", x"0308", x"03D4", x"0561", x"06F4", x"08A0", x"09B1", x"093D", x"084D", x"07CE", x"075F", x"0755", x"07CC", x"06F5", x"0409", x"011C", x"FF31", x"FE4E", x"FF8B", x"025B", x"043B", x"04B0", x"04F7", x"04CC", x"040B", x"03CD", x"03DC", x"0323", x"0233", x"0173", x"0053", x"FF30", x"FED9", x"FEFE", x"FF55", x"000C", x"005C", x"0011", x"FFB4", x"FF6B", x"FEED", x"FEDC", x"FEF0", x"FE8F", x"FE0F", x"FDB6", x"FD27", x"FCE3", x"FD85", x"FE41", x"FEBD", x"FF22", x"FEB3", x"FD34", x"FC45", x"FC79", x"FD5D", x"FF57", x"01BE", x"0241", x"00F3", x"FF85", x"FE6C", x"FE10", x"FFD9", x"0284", x"03FF", x"0485", x"0470", x"02E1", x"008B", x"FEAA", x"FCB0", x"FAAA", x"FA00", x"FA4E", x"FB37", x"FD92", x"00DF", x"03AD", x"062C", x"0836", x"088F", x"07DE", x"0751", x"061E", x"0487", x"041A", x"045C", x"0433", x"0477", x"04DF", x"0464", x"042B", x"057A", x"06FC", x"0860", x"09DC", x"0A44", x"0956", x"08ED", x"0931", x"094C", x"09B9", x"0999", x"074E", x"03D7", x"012F", x"FF6F", x"FF6D", x"01F9", x"0516", x"0706", x"0871", x"093A", x"08D4", x"08B1", x"0954", x"0982", x"099C", x"0A41", x"0AA3", x"0ACE", x"0BFF", x"0D66", x"0E7E", x"103A", x"1224", x"1334", x"1420", x"1507", x"14C7", x"1421", x"140E", x"13C2", x"12E8", x"124A", x"1153", x"0FF3", x"0F83", x"0FF3", x"1038", x"107C", x"1024", x"0E5E", x"0C64", x"0B66", x"0B20", x"0C26", x"0E98", x"1012", x"0F52", x"0DC8", x"0BC1", x"09D4", x"0A55", x"0CFE", x"0ED9", x"0F7A", x"0F69", x"0D7A", x"0A72", x"0835", x"05EC", x"0272", x"FF71", x"FD3F", x"FB07", x"FA18", x"FB0B", x"FBFA", x"FCAE", x"FDF8", x"FE8E", x"FDDC", x"FD51", x"FCA6", x"FB4A", x"FAC2", x"FB88", x"FC48", x"FD04", x"FDF7", x"FDED", x"FD1B", x"FCE2", x"FCC2", x"FC71", x"FCA1", x"FCAB", x"FBD3", x"FB60", x"FBBB", x"FC38", x"FD77", x"FF52", x"FF80", x"FDE8", x"FC2E", x"FAC9", x"FA5E", x"FCC1", x"00D7", x"0415", x"0665", x"0806", x"07F2", x"06C7", x"05ED", x"0494", x"029F", x"013A", x"006A", x"FF8E", x"FF83", x"0064", x"015C", x"02A8", x"0460", x"057E", x"061F", x"06CD", x"06FA", x"0692", x"065E", x"05C2", x"0463", x"030E", x"019F", x"FFA5", x"FE08", x"FD2A", x"FC15", x"FB36", x"FAB5", x"F96C", x"F775", x"F670", x"F621", x"F683", x"F891", x"FB04", x"FB91", x"FACD", x"F9E2", x"F897", x"F871", x"FAF5", x"FE29", x"007B", x"0298", x"03C8", x"0312", x"01DE", x"00AF", x"FE51", x"FBC1", x"FA62", x"F977", x"F96A", x"FB71", x"FE7C", x"015D", x"0501", x"0886", x"0A94", x"0C17", x"0D71", x"0D48", x"0C9C", x"0D1A", x"0DE0", x"0E90", x"102A", x"1165", x"112F", x"1141", x"1219", x"12A1", x"1321", x"13B0", x"129D", x"1082", x"0F38", x"0E87", x"0E50", x"0F1A", x"0F4A", x"0D30", x"0A34", x"075B", x"050D", x"0518", x"07F6", x"0B7E", x"0E7E", x"1127", x"1234", x"11A5", x"1117", x"104B", x"0E7F", x"0CC6", x"0B1C", x"08B4", x"0687", x"0548", x"03BF", x"021B", x"014C", x"0045", x"FED0", x"FE1D", x"FD5B", x"FBA3", x"FA1D", x"F93C", x"F80A", x"F754", x"F776", x"F72C", x"F6CB", x"F76A", x"F858", x"F93F", x"FA9F", x"FB66", x"FADC", x"FA70", x"FA69", x"FAA8", x"FC6A", x"FF72", x"0151", x"01A8", x"0143", x"FF99", x"FE04", x"FF20", x"01C9", x"03E4", x"05A5", x"066E", x"04E8", x"02C6", x"016E", x"FF4B", x"FC44", x"F9DB", x"F778", x"F4EA", x"F430", x"F4DA", x"F526", x"F5B0", x"F6A8", x"F6B8", x"F650", x"F6A3", x"F69D", x"F605", x"F655", x"F733", x"F7E8", x"F920", x"FA94", x"FB1B", x"FB6D", x"FC0F", x"FC45", x"FC57", x"FCC3", x"FC9A", x"FBF4", x"FBDD", x"FBF7", x"FC04", x"FCFB", x"FDCD", x"FCDB", x"FAA2", x"F803", x"F507", x"F38C", x"F51B", x"F81E", x"FAFB", x"FDAC", x"FF3D", x"FED8", x"FDF7", x"FD30", x"FBB6", x"FA28", x"F93C", x"F848", x"F752", x"F733", x"F77D", x"F7DC", x"F8F2", x"FA51", x"FB31", x"FBFB", x"FC9F", x"FC77", x"FC0D", x"FBCF", x"FB14", x"FA2F", x"F9B2", x"F8FB", x"F802", x"F7C4", x"F7D3", x"F7BB", x"F854", x"F903", x"F8B3", x"F804", x"F7DB", x"F7AA", x"F87B", x"FB38", x"FDE4", x"FEF1", x"FEDB", x"FD97", x"FB4B", x"FAA0", x"FC83", x"FF12", x"01A9", x"0441", x"052B", x"0456", x"036C", x"0218", x"FFF6", x"FE3E", x"FD57", x"FC66", x"FC7D", x"FE28", x"0025", x"0255", x"053F", x"076A", x"084D", x"08E1", x"0873", x"065C", x"0426", x"0292", x"0114", x"00A3", x"01A1", x"023A", x"023B", x"029F", x"02E3", x"02CD", x"0378", x"0405", x"0340", x"0228", x"014E", x"0039", x"FFED", x"00A1", x"004F", x"FE3F", x"FB74", x"F7F1", x"F4EB", x"F4D6", x"F77D", x"FB02", x"FEFC", x"026E", x"03C8", x"03FB", x"045A", x"041C", x"037C", x"0351", x"02AF", x"0158", x"00BA", x"00B5", x"0087", x"00FB", x"020F", x"0288", x"0325", x"048E", x"0583", x"05D0", x"0644", x"060E", x"0519", x"04AF", x"04A2", x"0456", x"04B1", x"05CE", x"0695", x"07B4", x"092D", x"09C4", x"09C0", x"09FD", x"09D1", x"099B", x"0AFF", x"0CC9", x"0D57", x"0D0E", x"0B37", x"0730", x"037B", x"022B", x"01FB", x"0271", x"039F", x"036C", x"0123", x"FF0B", x"FD42", x"FADF", x"F8EA", x"F7AB", x"F5A1", x"F3E5", x"F3CB", x"F450", x"F516", x"F6EB", x"F878", x"F8DA", x"F914", x"F916", x"F7F8", x"F6DB", x"F64A", x"F592", x"F556", x"F641", x"F70C", x"F77E", x"F832", x"F82D", x"F730", x"F683", x"F5EB", x"F4CC", x"F442", x"F467", x"F419", x"F456", x"F626", x"F7AE", x"F844", x"F868", x"F731", x"F4CC", x"F41B", x"F609", x"F939", x"FD52", x"019E", x"03E5", x"0416", x"03B1", x"02B5", x"0139", x"00AB", x"00EA", x"013E", x"020F", x"0362", x"0477", x"05C9", x"0798", x"0937", x"0A89", x"0BB6", x"0C0A", x"0B50", x"0A67", x"08B1", x"0644", x"0411", x"01F2", x"FF95", x"FDC8", x"FC9D", x"FB13", x"F9BF", x"F93F", x"F893", x"F7AA", x"F793", x"F752", x"F6BF", x"F75B", x"F944", x"FA9B", x"FB5F", x"FB40", x"F8F5", x"F5D1", x"F470", x"F4D3", x"F64D", x"F90A", x"FBA8", x"FC69", x"FC47", x"FBED", x"FAB8", x"F94B", x"F863", x"F712", x"F569", x"F4D3", x"F4FE", x"F5BD", x"F7E6", x"FAB9", x"FCAE", x"FE41", x"FFAF", x"FFCC", x"FF4C", x"FF15", x"FE71", x"FD75", x"FDCD", x"FEBC", x"FF6E", x"00A0", x"0204", x"022D", x"0233", x"02B0", x"026B", x"01AB", x"01A2", x"0155", x"00EE", x"01FA", x"03C0", x"0447", x"03EB", x"0270", x"FF22", x"FC42", x"FC2B", x"FDEF", x"00BB", x"0461", x"06C7", x"06CC", x"0606", x"050D", x"0340", x"01AA", x"009E", x"FEBB", x"FC87", x"FB30", x"FA12", x"F955", x"F9D0", x"FAAC", x"FAE5", x"FB6B", x"FBD5", x"FB62", x"FAC3", x"FA30", x"F8CC", x"F751", x"F68A", x"F5AA", x"F536", x"F5D0", x"F67D", x"F6D2", x"F7AE", x"F84A", x"F7F2", x"F82F", x"F891", x"F7FC", x"F7FB", x"F986", x"FB01", x"FC7E", x"FE6B", x"FE78", x"FC50", x"FB04", x"FB30", x"FC04", x"FE95", x"0210", x"0345", x"02CC", x"023E", x"00A7", x"FE53", x"FCF8", x"FB82", x"F8E7", x"F718", x"F658", x"F59B", x"F60F", x"F7DE", x"F929", x"FA16", x"FBA0", x"FC7E", x"FCA1", x"FD60", x"FDCB", x"FD64", x"FDD1", x"FECA", x"FF35", x"0014", x"013E", x"00B5", x"FF56", x"FE67", x"FCD0", x"FB0B", x"FAEE", x"FADF", x"F9EB", x"FA28", x"FBB2", x"FC7F", x"FD4B", x"FDE0", x"FC0E", x"F8D1", x"F78D", x"F819", x"F9BF", x"FD23", x"00A3", x"01DA", x"01EE", x"01D3", x"00E4", x"FFB5", x"FF49", x"FEB0", x"FDA9", x"FD13", x"FC7A", x"FBEC", x"FC49", x"FD4C", x"FE60", x"FFC5", x"00DF", x"00F4", x"00E0", x"00B3", x"FF8A", x"FE23", x"FCE8", x"FB0C", x"F946", x"F8F6", x"F8F5", x"F86B", x"F874", x"F83D", x"F6B7", x"F591", x"F544", x"F428", x"F330", x"F40F", x"F594", x"F6F9", x"F919", x"FA0E", x"F85C", x"F64D", x"F5EB", x"F6A1", x"F93E", x"FD94", x"00EE", x"021C", x"026C", x"01B2", x"FFD2", x"FE79", x"FD57", x"FB63", x"F957", x"F814", x"F6F6", x"F71D", x"F947", x"FBD4", x"FDD7", x"FFCD", x"00C8", x"004F", x"0005", x"0001", x"FF5A", x"FF50", x"0099", x"0212", x"03EE", x"06D1", x"0900", x"09C4", x"0A69", x"0A97", x"098F", x"08D8", x"086E", x"06D5", x"050A", x"0457", x"036A", x"01ED", x"0096", x"FE27", x"FA07", x"F719", x"F69D", x"F7D5", x"FAFD", x"FFA3", x"031E", x"04FD", x"067E", x"0748", x"0712", x"0737", x"0761", x"06AD", x"05E2", x"056B", x"0498", x"041A", x"049F", x"0560", x"0653", x"0802", x"098C", x"0A99", x"0BA6", x"0C23", x"0BBC", x"0B4F", x"0AEE", x"0A52", x"0A9E", x"0BD3", x"0CB1", x"0D8D", x"0E71", x"0E12", x"0D20", x"0D0E", x"0CAD", x"0B5D", x"0B18", x"0B72", x"0B40", x"0BDB", x"0CDB", x"0B4E", x"07C5", x"0516", x"02CE", x"0151", x"0284", x"0495", x"04D8", x"049C", x"04A0", x"0365", x"01B4", x"00C9", x"FECD", x"FBB7", x"F9A5", x"F876", x"F79C", x"F881", x"FA84", x"FBD3", x"FCF6", x"FE1C", x"FE0B", x"FD61", x"FD12", x"FC16", x"FAD2", x"FA8E", x"FA84", x"FA7F", x"FBAD", x"FD03", x"FCFF", x"FCE4", x"FC92", x"FAE8", x"F9A5", x"F9DC", x"F95F", x"F873", x"F91C", x"FA28", x"FABB", x"FC45", x"FD5C", x"FB54", x"F889", x"F796", x"F7EC", x"FA20", x"FEDC", x"0324", x"04ED", x"05C0", x"05F1", x"04EF", x"0427", x"043A", x"0417", x"03FB", x"046E", x"04BF", x"04FD", x"05E9", x"06FD", x"0817", x"0970", x"0A04", x"09C3", x"096F", x"0897", x"0699", x"047D", x"01C7", x"FDEE", x"FAD1", x"F978", x"F87D", x"F828", x"F905", x"F92E", x"F85E", x"F8D2", x"F9B0", x"F93C", x"F922", x"FA07", x"FA63", x"FB22", x"FD42", x"FDC7", x"FB8F", x"F8FA", x"F6DF", x"F512", x"F583", x"F817", x"FA17", x"FB51", x"FCC5", x"FD97", x"FDBD", x"FE4F", x"FEC1", x"FE48", x"FDE9", x"FDCB", x"FDA7", x"FE8A", x"00CE", x"036A", x"0658", x"096F", x"0B86", x"0CCF", x"0E15", x"0EBF", x"0EB6", x"0EFA", x"0F64", x"0FA3", x"10FB", x"1330", x"14D0", x"15C8", x"163B", x"14E2", x"12A3", x"1138", x"101F", x"0EDF", x"0ECB", x"0F89", x"0FBC", x"1025", x"10AC", x"0F42", x"0C46", x"0A08", x"08D3", x"08CA", x"0AFE", x"0E5C", x"107F", x"11A9", x"123F", x"1172", x"0F80", x"0D85", x"0B3C", x"089D", x"06DD", x"05E7", x"0547", x"0560", x"0602", x"066A", x"06B6", x"06DC", x"064E", x"0550", x"0441", x"02BF", x"00EC", x"FF63", x"FD9C", x"FBF3", x"FB55", x"FB55", x"FB9C", x"FCA9", x"FDAC", x"FD84", x"FD58", x"FD9E", x"FD00", x"FC13", x"FC4D", x"FCB6", x"FD4A", x"FFBA", x"0276", x"02C3", x"01D0", x"0106", x"FFCD", x"FF8F", x"01D8", x"0451", x"050E", x"0593", x"05D1", x"049A", x"033D", x"023E", x"0026", x"FD71", x"FBC7", x"FABF", x"FA32", x"FB37", x"FD37", x"FF5C", x"01FE", x"04BA", x"068F", x"07BB", x"0832", x"07A5", x"06C9", x"05FF", x"04FF", x"046D", x"04DC", x"0524", x"053A", x"055F", x"0411", x"0143", x"FF24", x"FD9D", x"FBA6", x"FAFA", x"FBF8", x"FD04", x"FF0A", x"0300", x"05BB", x"0546", x"03AA", x"0171", x"FEC9", x"FE5E", x"00E0", x"033A", x"04AA", x"0627", x"0687", x"0566", x"0426", x"02B2", x"0060", x"FE70", x"FD86", x"FD2C", x"FD9E", x"FF07", x"00B4", x"029F", x"048A", x"05AA", x"064E", x"06CB", x"069A", x"060D", x"0592", x"041B", x"01C9", x"0069", x"FFEA", x"FFAB", x"00A4", x"01DE", x"0149", x"FFE7", x"FF83", x"FEC6", x"FDB8", x"FE04", x"FE8D", x"FE3F", x"FF30", x"0141", x"01B8", x"00AD", x"FFD4", x"FED7", x"FE5C", x"0071", x"0412", x"06EB", x"0929", x"0B14", x"0B95", x"0AEE", x"09CD", x"080F", x"05CE", x"03F1", x"02A9", x"01BE", x"0173", x"01A0", x"027F", x"0412", x"058A", x"0695", x"074A", x"0776", x"06F8", x"06B1", x"0669", x"0566", x"047E", x"047F", x"04DE", x"05DD", x"07EA", x"094F", x"08F3", x"0826", x"0711", x"050E", x"033D", x"0278", x"017C", x"0086", x"0101", x"0190", x"006E", x"FE65", x"FC51", x"FA0E", x"F94D", x"FB68", x"FEE8", x"023F", x"05B0", x"089C", x"0A02", x"0A4A", x"09EB", x"0894", x"06C6", x"0582", x"04BB", x"0433", x"041A", x"0462", x"0503", x"0620", x"079C", x"0913", x"0A6E", x"0B54", x"0BF0", x"0C90", x"0D47", x"0DF4", x"0EFA", x"1042", x"1139", x"1236", x"1348", x"135D", x"127F", x"11C8", x"10CD", x"0F3E", x"0E3B", x"0DEB", x"0D2B", x"0D0D", x"0E60", x"0F08", x"0D96", x"0B26", x"07D5", x"03DB", x"01AB", x"0243", x"035C", x"041E", x"0511", x"052E", x"03CC", x"0223", x"004C", x"FDA2", x"FB22", x"F9E0", x"F963", x"F971", x"FA41", x"FB4E", x"FC30", x"FD2A", x"FE03", x"FE8D", x"FEBD", x"FE85", x"FE28", x"FDDF", x"FD37", x"FC4D", x"FBD5", x"FB8F", x"FB8A", x"FC9E", x"FE0C", x"FE0A", x"FD5D", x"FCDE", x"FB91", x"FA0E", x"F9DD", x"F9E1", x"F947", x"FA68", x"FD4B", x"FF0E", x"FF9B", x"FFA4", x"FE2B", x"FC2D", x"FCF0", x"FFD1", x"0274", x"04FF", x"077F", x"0879", x"089A", x"091D", x"0950", x"08D3", x"08D0", x"0969", x"0A28", x"0B39", x"0CB2", x"0E1D", x"0FBD", x"1131", x"122C", x"129B", x"1215", x"1097", x"0EBD", x"0C83", x"0918", x"0579", x"0263", x"FFA2", x"FE24", x"FEDB", x"FFE3", x"FFC5", x"FF99", x"FEFA", x"FD0F", x"FB67", x"FAE5", x"F9E3", x"F900", x"FA28", x"FBFE", x"FC5E", x"FBD6", x"FA29", x"F6A2", x"F380", x"F30C", x"F439", x"F5EA", x"F862", x"FAB8", x"FBC4", x"FBEB", x"FB94", x"FA74", x"F92A", x"F87D", x"F868", x"F892", x"F8A1", x"F8A3", x"F931", x"FA64", x"FBE6", x"FDAF", x"FF47", x"FFE3", x"0008", x"006E", x"009D", x"0067", x"00D7", x"0199", x"026D", x"044A", x"0721", x"090D", x"09EF", x"0A9E", x"0A48", x"08D8", x"07EA", x"0726", x"0572", x"0450", x"04B8", x"0500", x"042A", x"02D9", x"006B", x"FCF4", x"FB0C", x"FBBF", x"FD7C", x"FF76", x"01A8", x"02D3", x"0257", x"0139", x"FFB7", x"FD8F", x"FBB2", x"FADD", x"FAB2", x"FAC9", x"FB25", x"FB82", x"FBF0", x"FCC1", x"FDE9", x"FF2B", x"001A", x"0062", x"FFE4", x"FEDA", x"FD0E", x"FAFA", x"F93F", x"F7EC", x"F755", x"F83A", x"FA22", x"FBCC", x"FD65", x"FEDC", x"FF23", x"FE9F", x"FE84", x"FE16", x"FD1B", x"FD9A", x"FFB9", x"0149", x"0211", x"0204", x"FFD9", x"FC7C", x"FB2F", x"FBFE", x"FD4F", x"FF44", x"0159", x"01C1", x"00FE", x"005F", x"FF10", x"FCD0", x"FAE4", x"F967", x"F807", x"F7A7", x"F88A", x"FA02", x"FC23", x"FED1", x"0121", x"02E1", x"0404", x"0453", x"0417", x"03A8", x"02A0", x"0144", x"0015", x"FEA2", x"FD5F", x"FD1C", x"FCB4", x"FB27", x"F96F", x"F78D", x"F4CA", x"F307", x"F31B", x"F34E", x"F3E9", x"F6DA", x"FAA7", x"FD45", x"FF2F", x"FF7E", x"FC8B", x"F914", x"F834", x"F92A", x"FB1E", x"FE7B", x"0160", x"0212", x"01CD", x"0138", x"FF9E", x"FDCA", x"FCE8", x"FC89", x"FC8E", x"FD2E", x"FDF9", x"FEB7", x"FF84", x"0029", x"006E", x"0071", x"FFC6", x"FED9", x"FE3E", x"FD73", x"FBE0", x"FA54", x"F87E", x"F626", x"F514", x"F5B3", x"F63A", x"F681", x"F745", x"F726", x"F617", x"F62F", x"F6CC", x"F633", x"F61F", x"F7D0", x"F960", x"FA4C", x"FB43", x"FA48", x"F6D8", x"F433", x"F3FB", x"F502", x"F740", x"FA9F", x"FCD8", x"FD4F", x"FD0A", x"FBFD", x"F9AB", x"F741", x"F586", x"F438", x"F385", x"F38A", x"F3D2", x"F493", x"F5F4", x"F7D2", x"F9ED", x"FBF9", x"FD46", x"FE01", x"FE68", x"FE44", x"FDBE", x"FDA3", x"FDA9", x"FDFD", x"FF80", x"01E5", x"03B4", x"04F3", x"0599", x"048F", x"0267", x"00A3", x"FEE2", x"FCCF", x"FC26", x"FD22", x"FDD3", x"FDC9", x"FD0D", x"FA51", x"F673", x"F491", x"F58E", x"F80D", x"FBF0", x"0046", x"031A", x"044E", x"04F5", x"04E0", x"03E6", x"0335", x"02F8", x"02C4", x"02E7", x"0361", x"03CA", x"0458", x"052D", x"05BD", x"0635", x"06AF", x"06F6", x"0766", x"0849", x"08ED", x"0933", x"098E", x"0982", x"092F", x"0990", x"0A2C", x"0A0C", x"09F8", x"09FB", x"08D4", x"075E", x"066B", x"045D", x"0169", x"0001", x"FF9E", x"FEC9", x"FE3E", x"FD37", x"F9AC", x"F5B9", x"F498", x"F548", x"F6DF", x"F9B6", x"FBA9", x"FAC8", x"F93C", x"F839", x"F698", x"F538", x"F509", x"F492", x"F3D7", x"F445", x"F52B", x"F5C2", x"F705", x"F890", x"F95C", x"FA49", x"FB9E", x"FC48", x"FC89", x"FC95", x"FB83", x"F97B", x"F76C", x"F4F1", x"F2AD", x"F1A3", x"F134", x"F0D1", x"F12D", x"F15B", x"F089", x"F00E", x"EFF8", x"EEBF", x"EDDD", x"EECF", x"F040", x"F1D2", x"F45A", x"F584", x"F42B", x"F2FF", x"F390", x"F4DC", x"F7A6", x"FBB8", x"FE54", x"FED8", x"FEC6", x"FDCB", x"FBB7", x"FA21", x"F91A", x"F7E5", x"F745", x"F763", x"F761", x"F7A6", x"F860", x"F89F", x"F87F", x"F865", x"F7CB", x"F707", x"F6EE", x"F67F", x"F55D", x"F437", x"F295", x"F04D", x"EF63", x"EFDE", x"F045", x"F12E", x"F2DA", x"F357", x"F33B", x"F43F", x"F4B6", x"F38E", x"F340", x"F40A", x"F43C", x"F4AC", x"F56B", x"F373", x"EF42", x"EC94", x"EBF8", x"ECB0", x"EFC7", x"F3D2", x"F5EB", x"F68A", x"F74B", x"F76C", x"F6FD", x"F77F", x"F87B", x"F935", x"FA82", x"FC42", x"FD74", x"FE74", x"FFC2", x"0115", x"028F", x"048B", x"0671", x"07F4", x"0946", x"0A06", x"0A4C", x"0A66", x"0A31", x"09DB", x"0A44", x"0B44", x"0C5F", x"0DE6", x"0F1E", x"0EDC", x"0D8F", x"0C05", x"0963", x"0667", x"04E6", x"04AD", x"04AB", x"0511", x"04DE", x"0239", x"FE6D", x"FC1E", x"FB64", x"FC4B", x"FEFB", x"0201", x"0367", x"03F0", x"042B", x"03AE", x"02F5", x"02BE", x"0220", x"0100", x"FFB6", x"FE14", x"FC4B", x"FB4A", x"FAED", x"FAD1", x"FB3A", x"FBCA", x"FBC2", x"FBC5", x"FBAC", x"FA8D", x"F909", x"F7C8", x"F65C", x"F56D", x"F61B", x"F723", x"F7C0", x"F8CC", x"F9A9", x"F927", x"F8D9", x"F906", x"F7CA", x"F657", x"F6BB", x"F7D5", x"F8F6", x"FB37", x"FC8B", x"FAE3", x"F8E5", x"F8B3", x"F937", x"FAF9", x"FE77", x"00CC", x"00DC", x"00CE", x"009F", x"FF49", x"FE4C", x"FDD7", x"FC74", x"FAF3", x"FAA9", x"FA65", x"FA35", x"FB0B", x"FBF9", x"FC5B", x"FD49", x"FE72", x"FEDA", x"FF14", x"FF05", x"FDE3", x"FC34", x"FAA4", x"F887", x"F68A", x"F54F", x"F431", x"F358", x"F33B", x"F2D3", x"F1E8", x"F1A3", x"F186", x"F0D7", x"F124", x"F2DA", x"F4A7", x"F715", x"FA35", x"FB68", x"FA88", x"F9B4", x"F962", x"F978", x"FB81", x"FE81", x"0025", x"00A0", x"00AF", x"FF85", x"FDE3", x"FD2C", x"FCA5", x"FC12", x"FC6D", x"FD28", x"FDB6", x"FEF2", x"009E", x"01B0", x"02BA", x"03F2", x"047A", x"04F9", x"060A", x"0698", x"0696", x"06AF", x"05F2", x"0458", x"0358", x"02B7", x"01C1", x"01B3", x"026A", x"024A", x"024B", x"0325", x"02FE", x"01C2", x"0183", x"01B4", x"0162", x"01DD", x"0235", x"FF93", x"FB65", x"F87E", x"F6FB", x"F75C", x"FABF", x"FEE6", x"010C", x"01FE", x"0252", x"0117", x"FF56", x"FE58", x"FD6D", x"FC87", x"FCDD", x"FE00", x"FF04", x"0078", x"0240", x"0391", x"04C9", x"0615", x"06C5", x"06CD", x"069A", x"05F3", x"051F", x"0482", x"03F0", x"0379", x"039F", x"0412", x"04A7", x"05A7", x"062F", x"0590", x"0495", x"035C", x"0142", x"FF22", x"FE4B", x"FDD6", x"FD92", x"FE07", x"FDAC", x"FB11", x"F836", x"F6DC", x"F70F", x"F98C", x"FE67", x"0319", x"060F", x"081C", x"0910", x"08AA", x"0833", x"0812", x"077F", x"0702", x"06FC", x"06DE", x"06E2", x"07BE", x"08B2", x"096B", x"0A75", x"0B37", x"0B7C", x"0C29", x"0D09", x"0D5C", x"0DC6", x"0E55", x"0E3C", x"0E4C", x"0F2B", x"0F9B", x"0FA7", x"102A", x"0FF5", x"0ED3", x"0E6D", x"0E22", x"0C81", x"0B0D", x"0A81", x"0973", x"089A", x"08E4", x"07E4", x"04BC", x"0231", x"00CA", x"FFED", x"00F9", x"0368", x"0430", x"034C", x"0253", x"0098", x"FE74", x"FD9D", x"FD6D", x"FCCE", x"FCBF", x"FD31", x"FD23", x"FD8C", x"FEE4", x"0023", x"0181", x"0398", x"0554", x"068D", x"07E6", x"089A", x"0827", x"0775", x"0634", x"03F8", x"01E2", x"0024", x"FE4E", x"FD50", x"FD86", x"FD8A", x"FDC9", x"FEC4", x"FEF0", x"FE1C", x"FDF3", x"FE29", x"FE6A", x"0046", x"031D", x"0460", x"047A", x"04CF", x"04E0", x"0579", x"0802", x"0AD5", x"0C26", x"0CB1", x"0C76", x"0AFD", x"09B1", x"095D", x"091E", x"091D", x"09BB", x"09F0", x"09B5", x"09F8", x"0A24", x"0A0A", x"0A52", x"0A9B", x"0A4A", x"0A31", x"0A68", x"0A20", x"09E9", x"09BC", x"08A1", x"06C6", x"051B", x"0314", x"0137", x"00D3", x"010E", x"0144", x"0265", x"03EF", x"0423", x"03DE", x"03CC", x"02F1", x"01F1", x"0229", x"01DA", x"FF62", x"FC52", x"F998", x"F750", x"F72E", x"F9C5", x"FC83", x"FE22", x"FF1B", x"FF13", x"FE28", x"FDF5", x"FEDE", x"0002", x"01B8", x"03E3", x"0584", x"06BE", x"0805", x"08E1", x"0950", x"09FD", x"0AA1", x"0B20", x"0C1B", x"0D67", x"0E63", x"0F58", x"0FFE", x"0FC8", x"0F48", x"0EE1", x"0E67", x"0E33", x"0EBC", x"0EEA", x"0E8D", x"0E62", x"0DC4", x"0C01", x"0A5C", x"093F", x"0806", x"07A6", x"088B", x"089E", x"06E4", x"04E6", x"0359", x"0255", x"038E", x"06C4", x"0991", x"0B45", x"0C84", x"0CB1", x"0BD5", x"0B35", x"0A93", x"0947", x"07CA", x"0626", x"03DA", x"0198", x"0018", x"FF2E", x"FEF9", x"FFB7", x"0073", x"00F4", x"0186", x"01C1", x"0185", x"0173", x"013C", x"00C7", x"00CC", x"015A", x"01DA", x"02F8", x"0454", x"04D8", x"050B", x"05C1", x"05C8", x"0504", x"04C2", x"042D", x"02F0", x"02E7", x"03CF", x"0346", x"01B1", x"0043", x"FE57", x"FD15", x"FE8A", x"0141", x"033C", x"04EF", x"05F2", x"0541", x"0456", x"0427", x"03A3", x"0301", x"02EC", x"024B", x"0142", x"015F", x"022D", x"0327", x"051F", x"075D", x"088F", x"0981", x"0A54", x"09C5", x"0864", x"070C", x"04D9", x"023B", x"0066", x"FEAA", x"FCA8", x"FBC4", x"FB64", x"FAA4", x"FAC3", x"FBA9", x"FB57", x"FA8B", x"FA34", x"F956", x"F8BF", x"FA94", x"FD28", x"FE6A", x"FF3E", x"FF9D", x"FEE4", x"FF09", x"012F", x"0355", x"049F", x"058C", x"056D", x"0404", x"0309", x"0280", x"01DD", x"01A1", x"0197", x"00E2", x"002D", x"FFEB", x"FFC9", x"002D", x"0152", x"0220", x"0291", x"032F", x"0371", x"0373", x"03E5", x"040A", x"033F", x"0267", x"0169", x"0008", x"FFCE", x"00EB", x"01DE", x"0302", x"050B", x"0641", x"0673", x"06CD", x"0656", x"0426", x"0296", x"0212", x"00A2", x"FE4D", x"FBEF", x"F88E", x"F550", x"F4FA", x"F713", x"F9B0", x"FC82", x"FEA0", x"FEA2", x"FDD0", x"FD93", x"FD83", x"FDDF", x"FF22", x"001A", x"0077", x"0134", x"022A", x"02CE", x"03CE", x"04B9", x"0498", x"0428", x"042D", x"0423", x"045B", x"0558", x"060D", x"062A", x"0687", x"06BC", x"0690", x"06FB", x"0791", x"0734", x"069C", x"0654", x"0548", x"03C9", x"02E7", x"01B1", x"FFFE", x"FF86", x"0011", x"FFA2", x"FE65", x"FD11", x"FB4D", x"FA41", x"FBF9", x"FF8B", x"030F", x"0634", x"0876", x"08ED", x"0855", x"07B4", x"0711", x"0693", x"069A", x"06BA", x"0672", x"05FE", x"0566", x"04DF", x"04CA", x"04CC", x"0496", x"0464", x"0425", x"0407", x"04B2", x"0613", x"0753", x"08AD", x"09F9", x"0A87", x"0AE3", x"0BBA", x"0BCB", x"0ACB", x"09F1", x"08F7", x"0722", x"05D5", x"0504", x"0300", x"00BE", x"FFEF", x"FF40", x"FD94", x"FC08", x"F9F4", x"F6D8", x"F512", x"F616", x"F7F5", x"FA0C", x"FC4E", x"FD24", x"FC5E", x"FBCF", x"FB9E", x"FB47", x"FBAF", x"FC5B", x"FC0E", x"FB98", x"FB82", x"FB41", x"FB58", x"FC61", x"FD0E", x"FD13", x"FD73", x"FD90", x"FCE0", x"FC7B", x"FBEB", x"FA33", x"F833", x"F656", x"F3A1", x"F10E", x"EF85", x"EDE2", x"EC40", x"EC06", x"EC25", x"EBB2", x"EC01", x"ECCF", x"ECE9", x"EE42", x"F1D0", x"F56F", x"F80F", x"FA42", x"FAE0", x"FA1D", x"FA9E", x"FCE1", x"FF26", x"0125", x"02AA", x"0279", x"013B", x"003D", x"FF7F", x"FEF7", x"FF09", x"FEF7", x"FE43", x"FD5D", x"FC45", x"FB1D", x"FAB9", x"FACA", x"FA72", x"FA27", x"F9DE", x"F933", x"F8EC", x"F959", x"F939", x"F85D", x"F74B", x"F554", x"F2F5", x"F206", x"F20B", x"F215", x"F31C", x"F4E8", x"F5E7", x"F6BD", x"F801", x"F7D5", x"F639", x"F56B", x"F4FD", x"F3BB", x"F264", x"F0E2", x"EDD2", x"EB1F", x"EB1C", x"ECE9", x"EF8C", x"F2DF", x"F554", x"F5D6", x"F5DE", x"F656", x"F6F0", x"F875", x"FAE2", x"FCFC", x"FE84", x"0013", x"0117", x"01CE", x"02FF", x"042A", x"04BF", x"05A4", x"06E2", x"07F9", x"0979", x"0B39", x"0BFD", x"0BD8", x"0B49", x"0A00", x"086D", x"07D9", x"0769", x"067C", x"05EB", x"0563", x"0403", x"02C5", x"0222", x"00AD", x"FF0E", x"FEF1", x"FF50", x"FF01", x"FEB6", x"FE11", x"FC30", x"FB20", x"FC87", x"FF0C", x"01B9", x"049E", x"0679", x"0670", x"05D8", x"0517", x"03B7", x"0232", x"00F7", x"FF54", x"FD51", x"FB7C", x"F9A6", x"F821", x"F768", x"F71B", x"F6CC", x"F6A5", x"F64B", x"F5BC", x"F59B", x"F5B7", x"F599", x"F5A1", x"F589", x"F4E2", x"F498", x"F513", x"F533", x"F51B", x"F586", x"F54D", x"F451", x"F407", x"F3C6", x"F254", x"F15D", x"F1EB", x"F216", x"F1F9", x"F239", x"F15B", x"EF5D", x"EF4E", x"F1AB", x"F4C3", x"F86D", x"FC15", x"FD6F", x"FCF5", x"FC58", x"FB61", x"F9E9", x"F903", x"F83F", x"F6E3", x"F5FE", x"F5C9", x"F5E2", x"F6D8", x"F8D1", x"FA84", x"FBF6", x"FD40", x"FD7D", x"FCEE", x"FC62", x"FB39", x"F95B", x"F7BC", x"F5D2", x"F352", x"F1A7", x"F0A4", x"EF27", x"EE06", x"EDC3", x"ECD7", x"EBD4", x"EC13", x"EC2B", x"EBC5", x"ED41", x"F0A2", x"F3D8", x"F749", x"FA7D", x"FB3D", x"FA6C", x"FB02", x"FC9B", x"FE0E", x"FFDD", x"0111", x"0024", x"FE76", x"FD68", x"FC62", x"FB63", x"FB1B", x"FAD4", x"FA3F", x"FA1A", x"FA44", x"FA9A", x"FB77", x"FCA3", x"FD9C", x"FE85", x"FF26", x"FF59", x"FFBA", x"0068", x"00A9", x"00C1", x"00C3", x"FFFE", x"FF65", x"FFF3", x"00C1", x"0135", x"01EA", x"022C", x"0125", x"005C", x"0015", x"FEA8", x"FCC4", x"FBE0", x"FB0B", x"F972", x"F81F", x"F614", x"F23B", x"EEC6", x"EDCD", x"EE50", x"EFCC", x"F24C", x"F3FF", x"F428", x"F437", x"F4C9", x"F544", x"F60C", x"F761", x"F86C", x"F93D", x"FA27", x"FADF", x"FB6E", x"FC3A", x"FCE8", x"FD4A", x"FDAC", x"FDC2", x"FDBA", x"FE52", x"FF30", x"FF9E", x"FFE1", x"FF9F", x"FE49", x"FCEA", x"FC25", x"FADF", x"F912", x"F793", x"F598", x"F2F5", x"F185", x"F0F0", x"EFEF", x"EFB7", x"F142", x"F2C0", x"F3B2", x"F4D2", x"F473", x"F223", x"F0DC", x"F1F2", x"F3F1", x"F6EA", x"FAA6", x"FCE6", x"FD72", x"FE26", x"FEF2", x"FF16", x"FFB2", x"00C6", x"014F", x"01AB", x"0245", x"025C", x"0207", x"0201", x"01CE", x"0162", x"0130", x"0103", x"00DF", x"0174", x"02A4", x"03F2", x"05B7", x"075E", x"084D", x"090E", x"09A5", x"0947", x"087F", x"07EF", x"06AA", x"052E", x"0492", x"03B4", x"01F8", x"00FE", x"00A7", x"FFB7", x"FEB8", x"FDD0", x"FB0F", x"F76A", x"F5B2", x"F5E3", x"F74F", x"FA77", x"FDE5", x"FF63", x"FFC9", x"0036", x"FFE7", x"FF29", x"FEDC", x"FE3D", x"FD1C", x"FC8E", x"FC8D", x"FCA5", x"FD66", x"FE91", x"FF61", x"0036", x"011B", x"0180", x"01D3", x"023D", x"01EB", x"0101", x"FFE7", x"FDEA", x"FB7A", x"F9BD", x"F822", x"F636", x"F50B", x"F418", x"F299", x"F223", x"F336", x"F432", x"F57E", x"F873", x"FB89", x"FDFD", x"00EC", x"02D2", x"01AC", x"FFC3", x"FF3D", x"FF61", x"00C0", x"03E6", x"065E", x"06A9", x"06C5", x"071B", x"06C8", x"0694", x"06E2", x"0650", x"0544", x"051D", x"055F", x"05AC", x"0660", x"070E", x"06FE", x"06A4", x"0610", x"0540", x"047F", x"040A", x"0377", x"02D5", x"01D6", x"001E", x"FEB1", x"FE13", x"FDEB", x"FE66", x"FF94", x"0003", x"FFAB", x"FFF1", x"0038", x"FF63", x"FEA6", x"FE23", x"FC8A", x"FAA3", x"F958", x"F6B0", x"F253", x"EEF1", x"ED79", x"ED61", x"EF89", x"F346", x"F5B4", x"F671", x"F738", x"F7D0", x"F80B", x"F8FD", x"FA87", x"FBB8", x"FD20", x"FF4B", x"015A", x"0355", x"0571", x"0786", x"0963", x"0B1F", x"0C50", x"0D08", x"0D87", x"0D94", x"0D5A", x"0D11", x"0C0C", x"0A5E", x"095E", x"08D7", x"0838", x"0808", x"080A", x"06C9", x"056C", x"055C", x"0551", x"04CE", x"0557", x"0653", x"0678", x"0737", x"0870", x"0791", x"052D", x"03D7", x"0372", x"03BD", x"05F7", x"08BF", x"0981", x"0936", x"0929", x"0881", x"075A", x"06CC", x"060B", x"04B9", x"03E1", x"039D", x"0309", x"025A", x"01A2", x"0077", x"FF21", x"FDE8", x"FC9E", x"FBD0", x"FBBF", x"FC07", x"FCE4", x"FE44", x"FF54", x"006B", x"0254", x"043E", x"059E", x"0719", x"07E3", x"0720", x"0694", x"06C3", x"0653", x"05BC", x"0627", x"0637", x"05AA", x"060D", x"0611", x"041E", x"01EF", x"013D", x"014A", x"02DC", x"066D", x"0945", x"09FA", x"09EF", x"096A", x"07F1", x"06BE", x"0609", x"04B8", x"034F", x"02DD", x"02EF", x"038E", x"051E", x"06B5", x"07D4", x"08A7", x"08F3", x"0886", x"0852", x"081D", x"0783", x"06D4", x"05D4", x"03C1", x"01BA", x"0054", x"FECE", x"FD76", x"FCAE", x"FB08", x"F8AE", x"F766", x"F702", x"F6DD", x"F85A", x"FB4F", x"FE13", x"011A", x"04E1", x"06BB", x"05FE", x"0498", x"02F5", x"0159", x"01E3", x"043D", x"05A8", x"05D8", x"05BB", x"04C3", x"0359", x"0326", x"0360", x"031B", x"030E", x"034F", x"0337", x"033F", x"03A4", x"03B5", x"039E", x"03A0", x"0369", x"034F", x"03E3", x"04B4", x"05D5", x"075B", x"0862", x"08B1", x"096C", x"0A44", x"0AB6", x"0B77", x"0BDF", x"0A5B", x"084E", x"0714", x"05DF", x"04DE", x"0566", x"05F7", x"056C", x"0565", x"056F", x"0320", x"FF4D", x"FBDA", x"F86A", x"F61E", x"F715", x"F9B5", x"FB62", x"FCC6", x"FE31", x"FE8B", x"FEC0", x"FFD7", x"0090", x"0074", x"00CC", x"016B", x"01B4", x"0233", x"030E", x"03CD", x"04C8", x"0646", x"07BD", x"092A", x"0A80", x"0B70", x"0C46", x"0CDF", x"0C9F", x"0C00", x"0BC2", x"0B61", x"0B00", x"0B01", x"0A04", x"0744", x"0488", x"0289", x"00D7", x"00A3", x"0261", x"041B", x"056C", x"0765", x"0884", x"074F", x"055E", x"03A3", x"01D0", x"019B", x"040A", x"06D5", x"08B2", x"0A79", x"0BBA", x"0C14", x"0CC8", x"0DCD", x"0E04", x"0D99", x"0D3E", x"0C6C", x"0B70", x"0AD2", x"0A31", x"099C", x"0960", x"0931", x"090C", x"09C8", x"0AF7", x"0C72", x"0EA4", x"10D2", x"11F7", x"1324", x"14BA", x"159C", x"1656", x"1738", x"1698", x"1464", x"129A", x"10D7", x"0E4B", x"0C7E", x"0B8B", x"09C5", x"0837", x"07F9", x"06C1", x"03CD", x"00F8", x"FE88", x"FC5C", x"FCE3", x"0003", x"02B6", x"0453", x"0587", x"0569", x"0432", x"03B7", x"0375", x"0243", x"011E", x"0082", x"FFCA", x"FF5F", x"FFD8", x"0057", x"00CD", x"0188", x"022B", x"023A", x"020B", x"0146", x"FFEB", x"FE7B", x"FCA2", x"FA75", x"F895", x"F727", x"F5DA", x"F545", x"F4FC", x"F3C0", x"F238", x"F153", x"F0AD", x"F0C7", x"F2A8", x"F533", x"F775", x"FA59", x"FD58", x"FE7F", x"FE4E", x"FD82", x"FBD7", x"FAA3", x"FC1A", x"FF32", x"020B", x"04A6", x"0637", x"05DC", x"04CF", x"0434", x"0338", x"01F8", x"013F", x"0090", x"FFBF", x"FF80", x"FF64", x"FED2", x"FE3C", x"FD6C", x"FC0E", x"FAEC", x"FA45", x"F9B1", x"F99F", x"FA15", x"F9EC", x"F989", x"FA06", x"FAD0", x"FBAD", x"FD4B", x"FE45", x"FD4B", x"FBED", x"FB14", x"F9E3", x"F966", x"FA65", x"FB03", x"FABB", x"FB09", x"FAD1", x"F862", x"F550", x"F2C8", x"F06E", x"F00C", x"F32E", x"F75E", x"FA93", x"FD7A", x"FF9B", x"0051", x"014A", x"0335", x"0482", x"054D", x"06B0", x"0834", x"0977", x"0B36", x"0D20", x"0E7C", x"0FAB", x"10EC", x"118F", x"11B3", x"1175", x"10C9", x"1017", x"0F6F", x"0EB2", x"0E31", x"0E39", x"0E64", x"0ECA", x"0F33", x"0E69", x"0C20", x"0971", x"06B4", x"042B", x"033B", x"0406", x"054D", x"0741", x"09C2", x"0B18", x"0A6E", x"08CD", x"0650", x"038D", x"028B", x"03B5", x"055A", x"06FC", x"0878", x"08C3", x"083D", x"0828", x"082F", x"07CB", x"076C", x"06BE", x"053A", x"0395", x"021B", x"0060", x"FED8", x"FDA0", x"FBF1", x"FA26", x"F8E7", x"F7D2", x"F6F7", x"F72D", x"F7B8", x"F819", x"F966", x"FB74", x"FCEB", x"FE0E", x"FECD", x"FDD2", x"FBBA", x"FA71", x"F975", x"F890", x"F903", x"FA65", x"FB61", x"FD07", x"FF6D", x"0063", x"FFA1", x"FE6A", x"FC79", x"FA81", x"FAF8", x"FD65", x"FFA3", x"0177", x"02C6", x"0257", x"0115", x"00AA", x"0058", x"FF78", x"FF05", x"FECB", x"FE25", x"FDDE", x"FE3D", x"FE37", x"FDE8", x"FDCF", x"FD86", x"FCE4", x"FC79", x"FBCF", x"FA95", x"F916", x"F749", x"F510", x"F301", x"F157", x"EFE8", x"EEFA", x"EE28", x"ECCE", x"EB16", x"E97C", x"E81C", x"E7C2", x"E95D", x"EC37", x"EFEA", x"F478", x"F8A2", x"FB10", x"FC09", x"FBD4", x"FA6C", x"F97B", x"FA69", x"FC4A", x"FE4E", x"0055", x"0173", x"0149", x"013E", x"01D6", x"0250", x"02C9", x"0376", x"0388", x"033F", x"0359", x"036B", x"0346", x"0357", x"0369", x"0328", x"034C", x"03EA", x"0473", x"055F", x"0683", x"06DA", x"06D1", x"0713", x"0719", x"06F7", x"074E", x"06F3", x"051D", x"0318", x"012A", x"FEEB", x"FD78", x"FD80", x"FD7F", x"FD74", x"FE1A", x"FDD1", x"FB1E", x"F770", x"F331", x"EE9F", x"EC0D", x"ECEE", x"EF0A", x"F136", x"F3A1", x"F513", x"F514", x"F57D", x"F697", x"F710", x"F791", x"F8D8", x"F9F7", x"FAEA", x"FC5A", x"FD8E", x"FE0D", x"FEDD", x"0032", x"0190", x"032E", x"04D1", x"0598", x"05C5", x"059C", x"04E1", x"0408", x"037D", x"02AC", x"0166", x"FFF0", x"FD91", x"FA60", x"F773", x"F510", x"F2E2", x"F1E8", x"F23B", x"F306", x"F499", x"F717", x"F8BB", x"F8BE", x"F7ED", x"F65E", x"F49D", x"F4BC", x"F6F5", x"F9C3", x"FCBF", x"FFB1", x"0173", x"0241", x"0323", x"03B3", x"0396", x"037E", x"0350", x"02A7", x"021F", x"01CB", x"0132", x"00D5", x"00F6", x"00F2", x"015C", x"0265", x"0361", x"042E", x"0563", x"0610", x"0615", x"06BA", x"07D7", x"0862", x"08E0", x"0904", x"073D", x"0475", x"0224", x"FF97", x"FCDF", x"FB7C", x"FAE3", x"FA41", x"FB0C", x"FCD3", x"FD31", x"FC21", x"FA94", x"F7F3", x"F5A6", x"F622", x"F881", x"FAE2", x"FD6C", x"FF59", x"FF79", x"FF0F", x"FF64", x"FF31", x"FE7F", x"FE32", x"FDBA", x"FD08", x"FD7E", x"FEB3", x"FFAB", x"00D7", x"01ED", x"0213", x"01FE", x"0226", x"01A6", x"00B4", x"FFE6", x"FE6F", x"FC7A", x"FB58", x"FAAD", x"F9BB", x"F933", x"F884", x"F67D", x"F415", x"F218", x"EFD4", x"EE06", x"EE0E", x"EF43", x"F175", x"F56A", x"F99B", x"FBF7", x"FCC8", x"FC4E", x"FA60", x"F8E1", x"F972", x"FAF6", x"FCA6", x"FEC6", x"003C", x"0084", x"00E0", x"0179", x"018B", x"01AF", x"0211", x"020D", x"01D7", x"01F7", x"0197", x"00E4", x"0060", x"FF93", x"FEA1", x"FE59", x"FE69", x"FE29", x"FE4F", x"FE4D", x"FD53", x"FC86", x"FCD0", x"FD40", x"FE0E", x"FF68", x"FF74", x"FDB9", x"FBC5", x"F9AB", x"F6E0", x"F4F6", x"F426", x"F31D", x"F2D2", x"F400", x"F48E", x"F395", x"F1F4", x"EF24", x"EB67", x"E96F", x"EA00", x"EB60", x"ED9E", x"F0A1", x"F2CA", x"F438", x"F679", x"F8BE", x"FA6E", x"FC84", x"FEC2", x"005A", x"0227", x"0429", x"0542", x"05C4", x"0651", x"0643", x"0632", x"0713", x"07ED", x"0835", x"0891", x"0864", x"0745", x"06DD", x"078C", x"080A", x"0878", x"08BD", x"071F", x"03ED", x"00E9", x"FDB3", x"FA3C", x"F841", x"F7D7", x"F83B", x"FA74", x"FE5E", x"013F", x"0263", x"025C", x"00A6", x"FE38", x"FD9B", x"FECA", x"0050", x"024C", x"0446", x"04D3", x"04A9", x"04F2", x"0502", x"04CB", x"04FE", x"04ED", x"0417", x"0325", x"01F8", x"000D", x"FE2A", x"FC59", x"FA32", x"F8A2", x"F826", x"F81B", x"F8EE", x"FAC5", x"FC67", x"FDC5", x"FFD6", x"01FA", x"0386", x"0534", x"0651", x"0588", x"0434", x"031E", x"017D", x"0001", x"FFE7", x"002C", x"00BA", x"030F", x"05EB", x"071A", x"06FA", x"0565", x"01AB", x"FE0B", x"FD03", x"FD67", x"FE72", x"006C", x"01A4", x"0114", x"0088", x"008D", x"0004", x"FFA3", x"FFE2", x"FF8A", x"FF03", x"FF5C", x"FFA3", x"FF5F", x"FF62", x"FF2E", x"FE43", x"FE05", x"FE40", x"FDEC", x"FD8D", x"FD2A", x"FB8C", x"F98C", x"F887", x"F792", x"F696", x"F673", x"F5CD", x"F39F", x"F184", x"EFD4", x"ED9A", x"EC5E", x"ED1D", x"EE64", x"F0D3", x"F586", x"FA48", x"FD1F", x"FEA7", x"FE37", x"FB35", x"F88C", x"F7EE", x"F7F8", x"F893", x"FA64", x"FBA8", x"FBCC", x"FC6B", x"FD14", x"FCB1", x"FC61", x"FCB6", x"FCEA", x"FD8F", x"FEF1", x"FFDD", x"002B", x"0063", x"002B", x"FFC3", x"0022", x"00A4", x"0113", x"01F5", x"0265", x"01CE", x"016F", x"01C0", x"01F0", x"02CC", x"044A", x"0432", x"02C6", x"0193", x"FFF7", x"FDB8", x"FC95", x"FBE4", x"FA79", x"FA36", x"FBC3", x"FCA4", x"FC50", x"FB51", x"F80F", x"F344", x"F066", x"EFC6", x"F008", x"F1AF", x"F442", x"F59A", x"F668", x"F7F4", x"F933", x"F9F5", x"FB79", x"FD1F", x"FE47", x"FFDC", x"0155", x"01E5", x"026E", x"033E", x"03AC", x"04C1", x"06EF", x"08CB", x"0A6C", x"0C41", x"0CA2", x"0BA3", x"0B4D", x"0B52", x"0AF1", x"0B4F", x"0BCC", x"0A5C", x"083E", x"06F3", x"04FB", x"0271", x"0105", x"FFC2", x"FE80", x"FFD7", x"037A", x"06A3", x"0903", x"0A52", x"08DD", x"061E", x"0510", x"0549", x"05E1", x"07AA", x"097B", x"09B3", x"0982", x"0994", x"0903", x"085C", x"0872", x"0835", x"078D", x"0729", x"0663", x"051C", x"0444", x"036D", x"024C", x"01F8", x"0277", x"02E1", x"03FC", x"058E", x"0615", x"0649", x"076D", x"08A5", x"09B4", x"0B70", x"0C5D", x"0B4D", x"09E9", x"0878", x"060F", x"03CB", x"028B", x"0113", x"0033", x"01A1", x"03CC", x"0544", x"067E", x"064E", x"03D8", x"019E", x"0129", x"0166", x"028A", x"04B3", x"05CF", x"0552", x"0504", x"049B", x"0380", x"030B", x"0324", x"02B1", x"02A8", x"037E", x"03D9", x"03CC", x"03E5", x"0314", x"01A5", x"0120", x"00FF", x"0088", x"0081", x"001F", x"FE58", x"FC81", x"FB9C", x"FAA3", x"FA01", x"FA1B", x"F91F", x"F6A2", x"F460", x"F1E6", x"EEEF", x"ED43", x"ECE2", x"ECBD", x"EE5F", x"F29E", x"F734", x"FB69", x"FF38", x"006E", x"FECC", x"FD48", x"FCC3", x"FC45", x"FD18", x"FF05", x"FFC8", x"FFCF", x"00A5", x"0118", x"00A0", x"00B0", x"00C9", x"0027", x"0009", x"0081", x"001C", x"FF4D", x"FEAC", x"FD93", x"FCA6", x"FCCA", x"FD0C", x"FCF4", x"FD32", x"FCF7", x"FC32", x"FC64", x"FDA0", x"FF05", x"0119", x"0337", x"036E", x"0274", x"014F", x"FF4E", x"FCE2", x"FB89", x"FA2A", x"F885", x"F8DB", x"FB21", x"FD55", x"FF83", x"00CC", x"FEC2", x"FAA3", x"F7D8", x"F673", x"F667", x"F909", x"FCAC", x"FF17", x"0135", x"03C5", x"052A", x"0602", x"0778", x"0878", x"08F2", x"0A12", x"0B15", x"0B49", x"0B97", x"0C05", x"0BE1", x"0C4B", x"0D4C", x"0DBF", x"0E27", x"0ECC", x"0E54", x"0D6D", x"0D9C", x"0DF6", x"0E4E", x"0F82", x"1007", x"0E6A", x"0C5B", x"0A57", x"0759", x"04CA", x"03A4", x"022E", x"0162", x"0397", x"0779", x"0B42", x"0F54", x"1190", x"0FD5", x"0CD1", x"0AFD", x"0997", x"0968", x"0B6E", x"0D07", x"0D1D", x"0DB0", x"0E52", x"0DDE", x"0D9F", x"0DE2", x"0D03", x"0BE1", x"0B61", x"0A05", x"07D5", x"05EE", x"0385", x"00AF", x"FF1D", x"FE5B", x"FD95", x"FDA4", x"FE0F", x"FD72", x"FD19", x"FDFE", x"FEF2", x"005F", x"02B4", x"03FB", x"0383", x"0307", x"01EB", x"FFE7", x"FEAA", x"FE31", x"FD36", x"FD67", x"FFEB", x"02CF", x"05B4", x"08B7", x"0911", x"0647", x"0351", x"0116", x"FF59", x"FFCB", x"0220", x"0389", x"043C", x"0555", x"055E", x"045D", x"03C9", x"030E", x"01AA", x"0123", x"014D", x"00DE", x"007C", x"0039", x"FF11", x"FDF8", x"FDC4", x"FD4C", x"FC9B", x"FC48", x"FB08", x"F8C2", x"F769", x"F6CF", x"F670", x"F747", x"F868", x"F78E", x"F5B6", x"F3FC", x"F19B", x"EFC8", x"F00F", x"F0B0", x"F114", x"F37A", x"F77E", x"FB9E", x"00AC", x"056E", x"0672", x"04BB", x"0324", x"0187", x"00AC", x"029A", x"056F", x"06B8", x"07DC", x"0931", x"0921", x"08B8", x"0937", x"0961", x"095F", x"0A99", x"0BDD", x"0C1C", x"0C27", x"0BCD", x"0A6E", x"0992", x"0972", x"08F6", x"088E", x"0874", x"0778", x"0651", x"066F", x"072D", x"0840", x"0A55", x"0BD5", x"0B62", x"0A40", x"08CE", x"064E", x"0419", x"028C", x"0002", x"FD34", x"FC06", x"FBF8", x"FC87", x"FE76", x"FF90", x"FDA1", x"FA47", x"F731", x"F43D", x"F316", x"F494", x"F6A1", x"F7F6", x"F9B8", x"FB1D", x"FB90", x"FC65", x"FDB9", x"FE8F", x"FFA8", x"014A", x"026C", x"0360", x"04D9", x"05CB", x"0671", x"07A2", x"087A", x"08A0", x"0910", x"0913", x"0798", x"063F", x"0595", x"04CE", x"04B0", x"057E", x"04E7", x"0288", x"FFF9", x"FCB7", x"F8E0", x"F670", x"F4F1", x"F2FE", x"F260", x"F408", x"F69C", x"FA60", x"FF6A", x"0270", x"0252", x"0145", x"FFDC", x"FE28", x"FEA0", x"011E", x"02CC", x"03EE", x"0570", x"05E7", x"0576", x"05E7", x"0642", x"05CC", x"061B", x"070E", x"0724", x"0725", x"073A", x"0621", x"04BA", x"046D", x"045D", x"0448", x"0500", x"0554", x"04A6", x"0498", x"055D", x"0638", x"07A0", x"092E", x"0916", x"07B6", x"05EE", x"0341", x"007D", x"FED7", x"FD5D", x"FBDF", x"FBB3", x"FCA2", x"FE0F", x"0126", x"04DB", x"0657", x"05D8", x"0493", x"022A", x"004B", x"012A", x"0335", x"0481", x"05F5", x"0721", x"06DE", x"06C2", x"0795", x"07ED", x"0813", x"092C", x"0A05", x"0A25", x"0AA6", x"0AB9", x"09D8", x"0951", x"0927", x"083B", x"0740", x"0628", x"03C0", x"00F3", x"FF31", x"FDC6", x"FD0B", x"FD99", x"FDA6", x"FBEB", x"F98E", x"F64D", x"F211", x"EF02", x"EDC5", x"EC8E", x"EC34", x"EDF0", x"F060", x"F3EB", x"F9CE", x"FF36", x"0125", x"00E1", x"FF33", x"FBE9", x"FA11", x"FB58", x"FD30", x"FE73", x"0059", x"01DA", x"0221", x"02F7", x"0462", x"04E9", x"0551", x"0649", x"0689", x"061A", x"05E4", x"0576", x"04F5", x"053D", x"05AB", x"0583", x"0554", x"04C9", x"03AA", x"0330", x"0393", x"0429", x"0587", x"0744", x"07B6", x"06B6", x"04D0", x"0149", x"FCDE", x"F979", x"F67B", x"F331", x"F0F0", x"EFC8", x"EEF8", x"EFEE", x"F2ED", x"F4EB", x"F4CA", x"F38F", x"F0CE", x"ED84", x"EC94", x"EE2E", x"F03A", x"F2DD", x"F5F3", x"F7F3", x"F939", x"FAF0", x"FC58", x"FD2F", x"FE79", x"FF8C", x"FFDF", x"007E", x"0162", x"0225", x"038B", x"058E", x"06C8", x"07AE", x"08B8", x"08C3", x"0803", x"07ED", x"07EC", x"07CE", x"08CB", x"09FC", x"0974", x"07D5", x"057A", x"01A8", x"FDBD", x"FB3B", x"F901", x"F6BD", x"F60C", x"F673", x"F7A6", x"FB29", x"0036", x"03CC", x"0595", x"0616", x"04A5", x"02A0", x"02A1", x"03D0", x"04DF", x"0651", x"07A7", x"077E", x"06D0", x"0657", x"0559", x"041C", x"0392", x"02D6", x"0199", x"0097", x"FF7E", x"FE41", x"FDC5", x"FDD9", x"FDBF", x"FDEE", x"FE52", x"FE1D", x"FE17", x"FF03", x"005E", x"0254", x"0501", x"0705", x"076B", x"06F4", x"0542", x"0276", x"0037", x"FEA2", x"FCE5", x"FBBA", x"FB8C", x"FB4B", x"FBF6", x"FEC7", x"01B3", x"0326", x"0383", x"0213", x"FEC6", x"FC98", x"FD14", x"FE79", x"0054", x"0299", x"0364", x"0265", x"0183", x"00A1", x"FF37", x"FE81", x"FE8E", x"FE37", x"FE0F", x"FE85", x"FE8C", x"FE5D", x"FEA3", x"FE5F", x"FD37", x"FC20", x"FA95", x"F84E", x"F6B5", x"F63B", x"F62B", x"F71C", x"F8B5", x"F913", x"F80C", x"F650", x"F369", x"F027", x"EE46", x"ED49", x"EC82", x"ECC2", x"ED9F", x"EE31", x"EFE3", x"F33E", x"F606", x"F754", x"F78E", x"F5B8", x"F28D", x"F0F0", x"F179", x"F291", x"F456", x"F687", x"F7A6", x"F7F7", x"F8C8", x"F99A", x"FA3F", x"FB83", x"FD05", x"FE08", x"FEE1", x"FF82", x"FFBA", x"000B", x"0094", x"008D", x"0035", x"FFB2", x"FE9D", x"FDA0", x"FDAE", x"FE69", x"FFE5", x"0279", x"051A", x"0691", x"072D", x"0677", x"03DF", x"00B3", x"FDD9", x"FA98", x"F79D", x"F5A1", x"F3AD", x"F1F9", x"F23B", x"F3DC", x"F4F0", x"F57B", x"F4CD", x"F1AE", x"EDE8", x"EC18", x"EBD3", x"EC91", x"EEE5", x"F1B4", x"F393", x"F56B", x"F798", x"F908", x"FA20", x"FBA7", x"FCE4", x"FDBF", x"FF10", x"005E", x"0169", x"02DA", x"0471", x"054B", x"05E1", x"064B", x"05E3", x"055D", x"05BE", x"069A", x"07FE", x"0A10", x"0B80", x"0B4E", x"09E6", x"0769", x"03F5", x"00D3", x"FE74", x"FC3B", x"FAA3", x"F9EC", x"F960", x"F99B", x"FBC5", x"FEA2", x"00E2", x"0253", x"0212", x"FF64", x"FCA1", x"FB73", x"FB0B", x"FB28", x"FC28", x"FCB2", x"FC37", x"FC1A", x"FC87", x"FCA3", x"FD1C", x"FE39", x"FEEC", x"FF12", x"FF16", x"FE73", x"FD73", x"FCE9", x"FCCB", x"FCB8", x"FD20", x"FD90", x"FDA9", x"FE10", x"FF18", x"0049", x"0215", x"040B", x"051D", x"051B", x"0474", x"02B8", x"0097", x"FF41", x"FE42", x"FD46", x"FD22", x"FD2C", x"FCB1", x"FD68", x"0026", x"030F", x"058D", x"076A", x"06AE", x"0372", x"00E6", x"FFE8", x"FF27", x"FF36", x"001C", x"FFCA", x"FEC1", x"FE9C", x"FE99", x"FDF5", x"FDFE", x"FEAC", x"FEFF", x"FF9D", x"00A7", x"011A", x"0134", x"0162", x"0101", x"FFEA", x"FEB3", x"FCD7", x"FA92", x"F8D7", x"F7AF", x"F6DF", x"F710", x"F77A", x"F6F4", x"F5AA", x"F3A4", x"F063", x"ED41", x"EB6A", x"EA60", x"EA4B", x"EBBC", x"ED72", x"EEE6", x"F1A6", x"F587", x"F8B6", x"FB37", x"FC9B", x"FB43", x"F857", x"F69D", x"F5D9", x"F553", x"F5BB", x"F661", x"F5D7", x"F4F8", x"F4B0", x"F423", x"F394", x"F3E9", x"F4A9", x"F548", x"F60C", x"F687", x"F687", x"F6BF", x"F6EF", x"F6D2", x"F6CB", x"F6C0", x"F649", x"F642", x"F706", x"F7CD", x"F8FF", x"FB0F", x"FCB1", x"FD4A", x"FD68", x"FC79", x"FA3B", x"F84E", x"F70C", x"F595", x"F479", x"F411", x"F334", x"F2B0", x"F43B", x"F6E3", x"F979", x"FBF6", x"FD0C", x"FB61", x"F918", x"F814", x"F7DC", x"F88D", x"FABE", x"FCDE", x"FE06", x"FF5E", x"00B2", x"0125", x"016A", x"01F8", x"0214", x"020E", x"027F", x"02CA", x"0327", x"0433", x"0547", x"060B", x"06E5", x"0766", x"06E1", x"0657", x"061C", x"05E8", x"0682", x"082B", x"095B", x"095B", x"0870", x"0649", x"0348", x"00F4", x"FF64", x"FE12", x"FD8F", x"FDAE", x"FDC7", x"FEFA", x"01FA", x"05A5", x"0962", x"0CF5", x"0E8F", x"0DED", x"0D5F", x"0D9C", x"0E04", x"0F1C", x"107B", x"105B", x"0EE7", x"0D9F", x"0BFA", x"09B8", x"07F9", x"0676", x"0490", x"02F2", x"01BC", x"0011", x"FE43", x"FCD1", x"FB2F", x"F9C0", x"F958", x"F95F", x"F9B2", x"FACF", x"FC52", x"FDB2", x"FFA9", x"01C3", x"02D8", x"02EE", x"0218", x"FFDA", x"FD44", x"FB84", x"FA40", x"F9B4", x"FA58", x"FB07", x"FB49", x"FCA7", x"FF3D", x"01E8", x"0543", x"085A", x"08FE", x"07E0", x"0783", x"07B2", x"0812", x"09A8", x"0B1F", x"0AB7", x"09AB", x"0932", x"07FF", x"065A", x"0544", x"03E2", x"01F5", x"0090", x"FF7A", x"FDED", x"FC99", x"FB70", x"F9DA", x"F84F", x"F738", x"F601", x"F536", x"F56F", x"F5E0", x"F6AA", x"F828", x"F959", x"F96D", x"F8E3", x"F735", x"F429", x"F15E", x"EF85", x"EE29", x"EE16", x"EF65", x"F06A", x"F166", x"F3AB", x"F697", x"F96B", x"FCE0", x"FF6D", x"FF68", x"FEA3", x"FEFA", x"FFD0", x"0185", x"049C", x"073C", x"0831", x"0902", x"09CB", x"09D7", x"0A13", x"0B1F", x"0C09", x"0CC1", x"0D6F", x"0D4B", x"0C42", x"0B33", x"09D8", x"0859", x"0736", x"0612", x"04D7", x"048B", x"0517", x"05DF", x"0785", x"09DB", x"0B6D", x"0C15", x"0C1F", x"0A6B", x"0763", x"0491", x"01D9", x"FEE3", x"FCC0", x"FAF0", x"F870", x"F68A", x"F64A", x"F6AC", x"F7A0", x"F950", x"F99A", x"F7CE", x"F639", x"F598", x"F57F", x"F6F1", x"F9C7", x"FC0B", x"FDBA", x"000E", x"022A", x"03AA", x"0579", x"074E", x"085A", x"0951", x"0A0B", x"09D0", x"092F", x"088B", x"0763", x"0622", x"0557", x"0450", x"0322", x"02B9", x"0277", x"0213", x"02B0", x"03FB", x"04A9", x"04EF", x"04A0", x"02B3", x"000C", x"FE26", x"FC8D", x"FB4F", x"FB2B", x"FB1E", x"FA93", x"FAEF", x"FC7B", x"FE21", x"0062", x"02C8", x"0351", x"027F", x"0253", x"02C7", x"0378", x"054D", x"071F", x"0736", x"06C1", x"06D1", x"06AE", x"06B0", x"07AA", x"089B", x"090C", x"09AB", x"09EB", x"0952", x"0889", x"0798", x"061A", x"04DD", x"042C", x"037A", x"0368", x"0447", x"0500", x"05BD", x"0720", x"084F", x"08AB", x"08D8", x"0826", x"0601", x"03F1", x"0297", x"0161", x"00FE", x"018E", x"015D", x"009F", x"00DA", x"01B0", x"02F1", x"05B0", x"0856", x"08EA", x"08AA", x"090C", x"096C", x"0AA0", x"0D5D", x"0F87", x"0FF2", x"102A", x"1037", x"0F87", x"0F61", x"101B", x"109C", x"110F", x"11D1", x"11EA", x"1151", x"10D2", x"0FC0", x"0DFF", x"0C47", x"0A1D", x"0758", x"0540", x"03CA", x"022F", x"014E", x"0158", x"00EB", x"0000", x"FF25", x"FCF1", x"F9A1", x"F707", x"F548", x"F416", x"F497", x"F628", x"F6F6", x"F7C3", x"F97B", x"FB22", x"FD14", x"FFF6", x"01B9", x"0151", x"008D", x"002A", x"FFB0", x"0073", x"0277", x"03B2", x"03FE", x"0489", x"04C4", x"049D", x"055E", x"06E1", x"0886", x"0A9C", x"0CAA", x"0DB9", x"0E2D", x"0E42", x"0D9B", x"0CD5", x"0C50", x"0B59", x"0A69", x"0A69", x"0A5A", x"09EC", x"0A04", x"09ED", x"08CC", x"076A", x"05B2", x"0269", x"FE9E", x"FB6A", x"F853", x"F5A4", x"F47F", x"F3B5", x"F2AD", x"F2CD", x"F420", x"F5B1", x"F83E", x"FB3B", x"FC60", x"FBE9", x"FB79", x"FAF9", x"FABC", x"FC24", x"FE26", x"FF48", x"0051", x"01B2", x"0294", x"036A", x"04D6", x"05ED", x"06A5", x"07AB", x"087A", x"08F5", x"09EA", x"0B09", x"0BA8", x"0C8A", x"0D4A", x"0D52", x"0D73", x"0E24", x"0E2A", x"0DED", x"0E2C", x"0E16", x"0D4A", x"0C94", x"0B2B", x"0829", x"04F1", x"0224", x"FF60", x"FD8F", x"FD1D", x"FCB6", x"FC51", x"FD26", x"FEA7", x"00A2", x"03E5", x"073F", x"08D7", x"0991", x"0A75", x"0B0F", x"0C22", x"0E4E", x"0FBF", x"0F7B", x"0E91", x"0D41", x"0B64", x"0A20", x"09E2", x"09C0", x"09C0", x"09FA", x"09A8", x"08DF", x"084A", x"0796", x"06F5", x"06EC", x"0703", x"0738", x"083E", x"09DE", x"0B39", x"0CCA", x"0E56", x"0ED4", x"0E8B", x"0DCB", x"0BA1", x"084C", x"0514", x"01F7", x"FF20", x"FDD5", x"FD92", x"FD09", x"FCEA", x"FD88", x"FE35", x"FFC8", x"02E5", x"05B4", x"06FC", x"07D8", x"085C", x"0832", x"08E6", x"0A80", x"0B13", x"0A7E", x"0998", x"07ED", x"058C", x"03BA", x"026D", x"0128", x"0056", x"FFE5", x"FF16", x"FE4B", x"FDD1", x"FD56", x"FD15", x"FD1A", x"FCB2", x"FC45", x"FC8D", x"FD40", x"FE41", x"0004", x"01AD", x"0265", x"028D", x"0212", x"0019", x"FD7D", x"FAF6", x"F829", x"F58C", x"F42D", x"F312", x"F1AE", x"F0F2", x"F0B8", x"F087", x"F14D", x"F322", x"F437", x"F478", x"F539", x"F63C", x"F790", x"FA18", x"FD11", x"FEB4", x"FF66", x"FFBD", x"FF63", x"FE93", x"FE48", x"FE71", x"FECC", x"FFB4", x"00BD", x"0163", x"01A2", x"01B4", x"018C", x"018F", x"0191", x"015A", x"0191", x"0279", x"03C1", x"0591", x"07E3", x"09AB", x"0A92", x"0AF1", x"0A48", x"0858", x"0606", x"038D", x"0088", x"FDA4", x"FB41", x"F877", x"F595", x"F3C1", x"F2C4", x"F292", x"F3CC", x"F57D", x"F5D9", x"F558", x"F51B", x"F504", x"F5B2", x"F7FA", x"FA9F", x"FC58", x"FDC9", x"FF38", x"FFF1", x"0071", x"0147", x"020E", x"02B0", x"039D", x"0483", x"04EB", x"0548", x"05A4", x"0614", x"06B5", x"0772", x"07F6", x"08A0", x"0998", x"0A87", x"0BC1", x"0D59", x"0EC5", x"0FB5", x"1052", x"0FD7", x"0E21", x"0BEE", x"098D", x"06FC", x"04FB", x"0393", x"01DB", x"0039", x"FF35", x"FE87", x"FE4E", x"FF4D", x"002F", x"FFD3", x"FF14", x"FE9C", x"FE39", x"FEBF", x"0094", x"01EA", x"01F1", x"0194", x"00D4", x"FF6E", x"FE83", x"FE88", x"FEB1", x"FF0A", x"FFC8", x"FFF7", x"FF3F", x"FE40", x"FCF0", x"FB5A", x"FA2E", x"F975", x"F8FE", x"F963", x"FA9F", x"FC21", x"FE19", x"0076", x"0259", x"0393", x"0440", x"03D1", x"026E", x"0118", x"FFD4", x"FEB0", x"FE47", x"FE53", x"FDFE", x"FDF6", x"FE85", x"FF0F", x"0017", x"0201", x"031A", x"02BF", x"0242", x"01CE", x"0138", x"01D5", x"0380", x"0427", x"03F6", x"040C", x"03C5", x"02EB", x"02B4", x"02B4", x"020F", x"019E", x"01B7", x"0147", x"0077", x"FFD9", x"FED9", x"FD62", x"FC30", x"FAB2", x"F8CA", x"F739", x"F61E", x"F557", x"F579", x"F655", x"F6DB", x"F6EA", x"F654", x"F4AB", x"F28A", x"F0E1", x"EF5E", x"EE56", x"EE35", x"EE4C", x"EE36", x"EEF6", x"F021", x"F130", x"F316", x"F540", x"F5BD", x"F4D7", x"F40A", x"F2EC", x"F22E", x"F347", x"F4CD", x"F4C1", x"F43B", x"F3FD", x"F30C", x"F250", x"F2DD", x"F36F", x"F3C7", x"F543", x"F746", x"F8BA", x"FA25", x"FB66", x"FB72", x"FB42", x"FB69", x"FB6B", x"FB92", x"FC91", x"FD88", x"FE65", x"FFDE", x"0147", x"01E7", x"021A", x"0161", x"FF0A", x"FC59", x"F9E5", x"F763", x"F580", x"F4A9", x"F376", x"F223", x"F1F5", x"F249", x"F338", x"F5E7", x"F8C0", x"F983", x"F931", x"F8D8", x"F7EA", x"F7E9", x"FA03", x"FBCD", x"FBF9", x"FC37", x"FC83", x"FBF9", x"FC04", x"FCEC", x"FCEE", x"FC97", x"FD36", x"FDCF", x"FE0E", x"FEDF", x"FF90", x"FF8C", x"FFC6", x"0024", x"FFFE", x"0000", x"003A", x"FFDB", x"FF79", x"FFAA", x"FFC3", x"FFF0", x"00AA", x"00D5", x"0030", x"FFC9", x"FF3A", x"FE61", x"FE79", x"FF19", x"FF07", x"FF3F", x"002F", x"00BA", x"01FA", x"04C7", x"06C8", x"0701", x"0734", x"073B", x"06E7", x"087A", x"0B7F", x"0C9A", x"0BB5", x"0A20", x"06DF", x"02CA", x"003B", x"FE67", x"FC14", x"FAAE", x"FA2D", x"F935", x"F8A8", x"F904", x"F8CE", x"F84E", x"F884", x"F87D", x"F84D", x"F971", x"FAEB", x"FC00", x"FDA3", x"FF86", x"004F", x"00D5", x"00FF", x"FF53", x"FC8C", x"FA26", x"F784", x"F55A", x"F4FD", x"F546", x"F550", x"F681", x"F853", x"F9F6", x"FCDE", x"0106", x"038E", x"04CC", x"0602", x"0655", x"0687", x"08DA", x"0B6C", x"0B95", x"0A88", x"0898", x"04DD", x"0119", x"FECC", x"FC2E", x"F909", x"F6F7", x"F50B", x"F2CD", x"F179", x"F0C1", x"EF66", x"EE82", x"EE46", x"EDB1", x"ED89", x"EE85", x"EF5A", x"F056", x"F266", x"F493", x"F65C", x"F878", x"F9B6", x"F920", x"F818", x"F6D0", x"F4EC", x"F3D5", x"F3EE", x"F389", x"F330", x"F3A5", x"F37F", x"F35C", x"F53F", x"F778", x"F837", x"F8D9", x"F948", x"F88F", x"F96D", x"FD3E", x"00CA", x"02E4", x"04C4", x"0506", x"0386", x"0307", x"037E", x"02DB", x"0249", x"02AD", x"0270", x"0248", x"034C", x"03E4", x"036A", x"0340", x"02CD", x"01B8", x"01A7", x"028A", x"02F8", x"03C8", x"0528", x"05C9", x"061E", x"06B2", x"05D5", x"0361", x"0097", x"FD01", x"F8D9", x"F611", x"F427", x"F203", x"F0CC", x"F089", x"EFD8", x"F06F", x"F33E", x"F5AC", x"F69F", x"F754", x"F6B4", x"F505", x"F5CA", x"F905", x"FBA1", x"FD9B", x"FF59", x"FF16", x"FDC8", x"FDDC", x"FE21", x"FD5A", x"FCEE", x"FC97", x"FB44", x"FA2A", x"F9CC", x"F8D1", x"F7BC", x"F729", x"F61E", x"F511", x"F52B", x"F5BB", x"F661", x"F80B", x"F9CB", x"FAEB", x"FC70", x"FDF1", x"FE24", x"FDDD", x"FD63", x"FB9B", x"F99A", x"F8BF", x"F7A8", x"F672", x"F664", x"F628", x"F526", x"F5B9", x"F7A2", x"F886", x"F936", x"FA25", x"F985", x"F913", x"FBAB", x"FF6B", x"0218", x"0468", x"0561", x"038E", x"0187", x"0103", x"004E", x"FFA0", x"001D", x"001C", x"FF3F", x"FF0E", x"FEFB", x"FE16", x"FDA6", x"FD7A", x"FC73", x"FBD9", x"FC52", x"FCA2", x"FD3C", x"FEF2", x"0057", x"014A", x"02E2", x"03D7", x"032C", x"023A", x"00CE", x"FE63", x"FCAF", x"FC49", x"FBC9", x"FBFC", x"FD78", x"FE84", x"FF6F", x"0214", x"04E7", x"0691", x"084F", x"097F", x"08FB", x"0995", x"0CC5", x"1012", x"12BB", x"1546", x"15BC", x"13EF", x"128B", x"1196", x"0FA8", x"0DF0", x"0CBD", x"0AA9", x"0894", x"0785", x"0630", x"048E", x"038B", x"020E", x"FFD5", x"FE2C", x"FCD5", x"FB23", x"FA6A", x"FA9F", x"FAB4", x"FB34", x"FC3B", x"FBEE", x"FA9C", x"F92C", x"F6FF", x"F4A3", x"F3C3", x"F38D", x"F33D", x"F404", x"F4E9", x"F47D", x"F480", x"F5AE", x"F63E", x"F677", x"F74D", x"F6CF", x"F570", x"F68D", x"F9E8", x"FD49", x"0108", x"044E", x"04B4", x"03B3", x"03B8", x"03B4", x"034F", x"03FE", x"04AF", x"0484", x"04FB", x"0614", x"0686", x"06E8", x"0794", x"072B", x"065B", x"0621", x"05BB", x"0509", x"0513", x"04FE", x"0441", x"03CA", x"032C", x"0143", x"FF00", x"FCA7", x"F988", x"F6DA", x"F562", x"F417", x"F33A", x"F39C", x"F3E5", x"F3C5", x"F528", x"F76E", x"F91A", x"FACD", x"FBED", x"FABB", x"F901", x"F976", x"FB41", x"FD77", x"008A", x"02A7", x"0250", x"017A", x"013A", x"009D", x"0035", x"00BB", x"0102", x"00F9", x"01AA", x"0299", x"0350", x"048D", x"05D4", x"065F", x"06BE", x"0731", x"06FF", x"06EE", x"075B", x"078F", x"07B0", x"0849", x"085B", x"07A8", x"06DD", x"0593", x"03B0", x"0256", x"017A", x"009B", x"00A3", x"019F", x"023D", x"02FC", x"04C2", x"0653", x"0761", x"08D6", x"0980", x"08BF", x"08E8", x"0B20", x"0E08", x"1149", x"148B", x"154A", x"1354", x"10D7", x"0E5C", x"0BB6", x"0A47", x"0A06", x"099B", x"094C", x"099E", x"0997", x"0957", x"09BB", x"0A10", x"0A1C", x"0AB1", x"0BAF", x"0C44", x"0D22", x"0E54", x"0F02", x"0F72", x"0FDB", x"0F10", x"0CEA", x"0A0D", x"069C", x"02F9", x"004B", x"FE68", x"FCFB", x"FCB0", x"FD1F", x"FD98", x"FED6", x"0115", x"0331", x"0537", x"0752", x"0811", x"077C", x"07E5", x"0988", x"0B65", x"0DB8", x"0FAA", x"0F24", x"0CD4", x"0AB7", x"087D", x"062E", x"04F1", x"0432", x"02EF", x"01FF", x"01BF", x"010A", x"004A", x"000B", x"FF81", x"FEA8", x"FE55", x"FE1B", x"FD64", x"FD2A", x"FD82", x"FE18", x"FF33", x"00A4", x"0116", x"0056", x"FEC4", x"FC77", x"FA1E", x"F851", x"F6C6", x"F592", x"F517", x"F4A8", x"F41B", x"F475", x"F552", x"F613", x"F761", x"F8A8", x"F84F", x"F779", x"F833", x"FA20", x"FCE5", x"00F9", x"042D", x"04A2", x"03B9", x"02A1", x"00CA", x"FF37", x"FF0B", x"FF2A", x"FF4F", x"00B0", x"02B3", x"044F", x"0638", x"083E", x"0954", x"0A4E", x"0BC7", x"0D01", x"0DF4", x"0F5B", x"1061", x"10AA", x"10E0", x"104B", x"0E2E", x"0B13", x"075B", x"02F4", x"FF0C", x"FC02", x"F965", x"F793", x"F6CF", x"F60B", x"F593", x"F668", x"F7B2", x"F911", x"FB05", x"FC4E", x"FBA3", x"FAF0", x"FBC2", x"FD9D", x"00AD", x"0518", x"083F", x"0907", x"0912", x"08A8", x"0770", x"06C8", x"073F", x"0792", x"0813", x"096C", x"0A90", x"0B1F", x"0C00", x"0CBA", x"0CEE", x"0D89", x"0EA5", x"0F4D", x"1011", x"1117", x"11BA", x"1231", x"12D5", x"12E7", x"11D2", x"1035", x"0E00", x"0B81", x"0965", x"0783", x"05AF", x"044F", x"0346", x"0236", x"01D0", x"0218", x"024A", x"02B4", x"0371", x"02EF", x"015C", x"006B", x"008A", x"0195", x"0464", x"07BE", x"0910", x"0887", x"06F4", x"0437", x"0140", x"FFC2", x"FF38", x"FED8", x"FF8A", x"00DD", x"01C1", x"02D3", x"045D", x"054A", x"05F9", x"077E", x"0914", x"0A44", x"0BCB", x"0D3D", x"0DEE", x"0EAF", x"0F99", x"0F71", x"0DFD", x"0BBE", x"089F", x"0573", x"032F", x"01CF", x"013C", x"01A8", x"0279", x"0354", x"04C2", x"0650", x"0795", x"0926", x"0A9B", x"0A8E", x"09E3", x"0A18", x"0B31", x"0D73", x"1171", x"152B", x"1675", x"160E", x"1499", x"11AD", x"0E7D", x"0C42", x"0A07", x"079E", x"0623", x"0521", x"0381", x"01E4", x"006F", x"FE45", x"FC3D", x"FB4A", x"FAC4", x"FA25", x"FA23", x"FA6E", x"FAB2", x"FB46", x"FC0B", x"FBD8", x"FA6A", x"F857", x"F613", x"F424", x"F2BE", x"F1E6", x"F1B3", x"F1BE", x"F1AF", x"F1CF", x"F220", x"F20E", x"F22E", x"F332", x"F3B7", x"F307", x"F22C", x"F1E8", x"F226", x"F443", x"F83C", x"FB90", x"FD06", x"FD7B", x"FCA2", x"FAA2", x"F92D", x"F8CA", x"F84C", x"F86E", x"F9AE", x"FB11", x"FC5B", x"FE3B", x"FFFC", x"0108", x"026C", x"0423", x"057A", x"06D9", x"0874", x"0987", x"0A23", x"0AAC", x"0A57", x"08BE", x"063F", x"02FE", x"FF4B", x"FC1C", x"F977", x"F751", x"F61C", x"F573", x"F4B8", x"F47E", x"F4F1", x"F57B", x"F69B", x"F88A", x"F98B", x"F917", x"F8BE", x"F914", x"FA49", x"FD8D", x"0242", x"05D5", x"078B", x"07EF", x"0695", x"03DC", x"01BA", x"006F", x"FF9A", x"FFE0", x"011A", x"01F0", x"024F", x"0299", x"024C", x"01A6", x"0192", x"01E3", x"0225", x"02C8", x"03DA", x"04E8", x"0646", x"0809", x"0952", x"09B9", x"094E", x"0861", x"0767", x"06D3", x"0695", x"06BE", x"0714", x"0734", x"0736", x"077C", x"0770", x"0749", x"079B", x"07ED", x"0725", x"05E9", x"04B7", x"03B9", x"03CE", x"05E3", x"0861", x"09C2", x"09EF", x"087F", x"0555", x"0216", x"FFF8", x"FE8F", x"FE1F", x"FED9", x"FFAD", x"0004", x"0075", x"00BF", x"0054", x"0033", x"00D2", x"0196", x"0267", x"0393", x"0464", x"0487", x"04D8", x"0529", x"04B5", x"0358", x"013C", x"FEA9", x"FC42", x"FAA3", x"F9E3", x"F9FF", x"FA99", x"FB79", x"FCC6", x"FE78", x"000E", x"01CC", x"03E6", x"055E", x"056F", x"04E1", x"042D", x"03C0", x"04E5", x"07EC", x"0AEA", x"0C90", x"0CBF", x"0B28", x"07C0", x"0432", x"014D", x"FEA1", x"FC91", x"FB9D", x"FADA", x"F9D4", x"F8F1", x"F811", x"F6AA", x"F5A9", x"F572", x"F55E", x"F514", x"F54D", x"F5D7", x"F6B3", x"F866", x"FAAD", x"FC34", x"FC62", x"FBBD", x"FAAA", x"F973", x"F86D", x"F7FC", x"F7BD", x"F743", x"F6D0", x"F69B", x"F633", x"F591", x"F599", x"F63F", x"F678", x"F5F3", x"F550", x"F4AD", x"F4D0", x"F735", x"FB97", x"FFF8", x"0347", x"054C", x"053D", x"0394", x"01EC", x"00DA", x"002A", x"0077", x"01AF", x"02AD", x"032C", x"03A0", x"03C1", x"03BA", x"0465", x"05AC", x"06B6", x"0789", x"0835", x"085B", x"083F", x"0831", x"07AB", x"05FE", x"0326", x"FF91", x"FBC4", x"F870", x"F5FF", x"F4B8", x"F46F", x"F49F", x"F506", x"F5BC", x"F672", x"F71A", x"F85B", x"F9F9", x"FA8E", x"F9F7", x"F906", x"F7F5", x"F7A4", x"F964", x"FCA6", x"FFAB", x"01E2", x"030A", x"0251", x"0022", x"FDF1", x"FC08", x"FAB0", x"FA97", x"FB61", x"FBF0", x"FC49", x"FC6A", x"FC23", x"FBD4", x"FC4A", x"FCF7", x"FD68", x"FDCD", x"FDE6", x"FD7B", x"FD2B", x"FD44", x"FCFD", x"FBF1", x"FA37", x"F7D4", x"F54B", x"F344", x"F217", x"F196", x"F18D", x"F1B0", x"F1F3", x"F284", x"F330", x"F42A", x"F59B", x"F6EB", x"F73E", x"F6DD", x"F666", x"F63A", x"F76D", x"FA7A", x"FE4F", x"0164", x"0337", x"0321", x"00F8", x"FDEB", x"FB31", x"F90D", x"F81F", x"F890", x"F9AE", x"FAC2", x"FC0E", x"FD28", x"FDC4", x"FEA0", x"FFFC", x"0149", x"0265", x"038B", x"0428", x"0444", x"0495", x"0525", x"04EF", x"03B4", x"019D", x"FEF3", x"FC4C", x"FAA4", x"FA3C", x"FABB", x"FBAD", x"FCE1", x"FE4D", x"FFB6", x"0106", x"02C9", x"04F1", x"069A", x"0756", x"0770", x"0727", x"071C", x"08DC", x"0C94", x"108E", x"13DD", x"15B3", x"153F", x"1292", x"0F4F", x"0C12", x"08C6", x"064B", x"04B6", x"02FF", x"010E", x"FF5E", x"FD61", x"FB14", x"F9B7", x"F944", x"F8BE", x"F844", x"F7DD", x"F6DF", x"F5BB", x"F5A0", x"F60D", x"F604", x"F55E", x"F41F", x"F214", x"EFF8", x"EE6F", x"ED8F", x"ED21", x"ED04", x"ED20", x"ED63", x"EDC0", x"EE35", x"EF76", x"F18E", x"F36A", x"F4AE", x"F5BC", x"F6B0", x"F80E", x"FB7A", x"0080", x"054F", x"090C", x"0B5F", x"0B34", x"08E6", x"05F6", x"02DB", x"FFB5", x"FDC0", x"FD1B", x"FCB9", x"FC84", x"FCB3", x"FCA9", x"FCB5", x"FDB2", x"FF51", x"00B6", x"01FB", x"02F7", x"034E", x"0370", x"03DB", x"03CD", x"02B5", x"0069", x"FD23", x"F942", x"F56E", x"F220", x"EFDC", x"EE6F", x"ED6F", x"ECE2", x"ECD6", x"ECB4", x"ECCD", x"EE24", x"F006", x"F143", x"F20E", x"F2BF", x"F30C", x"F465", x"F7F7", x"FC7E", x"007A", x"03B4", x"055F", x"04CF", x"0339", x"01B8", x"0023", x"FF29", x"FF6A", x"FFF9", x"0050", x"00D3", x"0111", x"00BA", x"00D0", x"016D", x"01F6", x"0295", x"0379", x"03C6", x"03C0", x"041E", x"049E", x"04BE", x"0484", x"0385", x"0186", x"FF4E", x"FD8A", x"FC5D", x"FC2E", x"FCB9", x"FD1A", x"FD61", x"FDA4", x"FDC5", x"FE60", x"0027", x"0229", x"0355", x"03D7", x"03BB", x"0330", x"03BC", x"0607", x"08ED", x"0B6F", x"0D0F", x"0CCA", x"0A8C", x"0766", x"0437", x"0160", x"FFAB", x"FF18", x"FEEC", x"FEE7", x"FF1C", x"FF17", x"FF32", x"FFF1", x"0137", x"0298", x"041D", x"0562", x"05EC", x"05FE", x"05FF", x"05D5", x"051F", x"039B", x"011B", x"FE00", x"FA98", x"F78D", x"F58C", x"F493", x"F441", x"F4A8", x"F5C2", x"F69E", x"F732", x"F872", x"FA0A", x"FB4A", x"FC48", x"FCEB", x"FC86", x"FC4D", x"FDF0", x"0153", x"057A", x"0A15", x"0DA8", x"0EDD", x"0E3F", x"0CC6", x"0A78", x"07FD", x"063A", x"04AD", x"02CD", x"0128", x"FF8B", x"FD57", x"FB3A", x"F9BC", x"F883", x"F75B", x"F6A0", x"F5E0", x"F4B8", x"F3E4", x"F3ED", x"F463", x"F4EB", x"F544", x"F53B", x"F4C5", x"F43C", x"F3F0", x"F403", x"F42B", x"F431", x"F44F", x"F45B", x"F3DB", x"F333", x"F338", x"F39D", x"F3B3", x"F3C1", x"F381", x"F2CE", x"F2E2", x"F510", x"F8BC", x"FCB0", x"0072", x"0304", x"0372", x"0277", x"00F5", x"FF1A", x"FD72", x"FCD5", x"FD10", x"FD90", x"FE66", x"FF8A", x"00CF", x"028F", x"052A", x"0811", x"0A85", x"0C3F", x"0D33", x"0D6D", x"0D47", x"0D2F", x"0CA7", x"0B02", x"07F2", x"0430", x"FFE8", x"FB6D", x"F7C0", x"F558", x"F3AE", x"F2C6", x"F302", x"F388", x"F38E", x"F428", x"F5DF", x"F7C7", x"F981", x"FB28", x"FBEB", x"FBD2", x"FCD7", x"FFD0", x"03BE", x"081D", x"0C4E", x"0EF0", x"0F96", x"0F34", x"0E1B", x"0C98", x"0B82", x"0B3F", x"0B43", x"0B6C", x"0BB9", x"0BC5", x"0BDE", x"0C6B", x"0D48", x"0E1D", x"0ECA", x"0ED5", x"0E3B", x"0D28", x"0C24", x"0B10", x"0A1F", x"08CE", x"06E1", x"04A3", x"0223", x"FFB1", x"FDFC", x"FD59", x"FD51", x"FDA1", x"FE49", x"FE55", x"FDAA", x"FD47", x"FD91", x"FDEF", x"FE30", x"FE3C", x"FD77", x"FC3A", x"FC09", x"FD25", x"FF08", x"012C", x"030A", x"03A0", x"02B5", x"00E2", x"FEB6", x"FCD2", x"FBEE", x"FC60", x"FDD1", x"FFDA", x"0233", x"04BF", x"0774", x"0A3A", x"0CF3", x"0F29", x"1081", x"10F8", x"10A0", x"0FAB", x"0E54", x"0CFF", x"0B15", x"087C", x"0589", x"0279", x"FF53", x"FCD2", x"FB86", x"FB04", x"FB44", x"FCB2", x"FEAF", x"0054", x"01FA", x"03FC", x"0606", x"07CB", x"0996", x"0A99", x"0A92", x"0A94", x"0BC9", x"0E2B", x"1160", x"14F3", x"1792", x"1860", x"1766", x"1533", x"1202", x"0E8F", x"0B76", x"08BC", x"0619", x"03A1", x"0148", x"FEED", x"FCFC", x"FBBC", x"FAF5", x"FA43", x"F9A1", x"F8F7", x"F839", x"F7EA", x"F874", x"F974", x"FA0D", x"FA2A", x"F9A5", x"F894", x"F74E", x"F690", x"F627", x"F5C6", x"F570", x"F572", x"F548", x"F4A0", x"F412", x"F414", x"F449", x"F49E", x"F519", x"F52B", x"F4A3", x"F4C7", x"F6C9", x"FA01", x"FDDE", x"01EF", x"050B", x"0631", x"05F6", x"04FD", x"030E", x"00EE", x"FFB5", x"FF3A", x"FF19", x"FFA4", x"00AD", x"01B8", x"0336", x"0598", x"0813", x"0A01", x"0B67", x"0BEF", x"0B8C", x"0B08", x"0AC5", x"0A31", x"0896", x"061D", x"02AD", x"FE83", x"FA33", x"F6B3", x"F3FE", x"F1F4", x"F0E0", x"F0C6", x"F0BE", x"F069", x"F0A0", x"F1AD", x"F2FC", x"F4A3", x"F691", x"F7AD", x"F83A", x"F9C9", x"FCEA", x"009C", x"04AB", x"08A3", x"0B2D", x"0C02", x"0BF9", x"0B08", x"091B", x"0737", x"0605", x"053B", x"04C5", x"04BB", x"04A6", x"048B", x"04E3", x"05E5", x"0718", x"085F", x"0985", x"0A85", x"0B7C", x"0CB3", x"0E17", x"0F26", x"0F3F", x"0E59", x"0CBE", x"0A82", x"080F", x"063B", x"0502", x"0406", x"03A7", x"03CA", x"033D", x"0229", x"01C3", x"021D", x"02AC", x"03C9", x"04CC", x"0463", x"0351", x"034A", x"0460", x"05F2", x"084F", x"0A8E", x"0B6D", x"0B21", x"0A4B", x"08AA", x"0656", x"0489", x"0358", x"0298", x"0282", x"0311", x"03F3", x"051A", x"06E1", x"08D8", x"0A6C", x"0B65", x"0BA8", x"0B20", x"0A3D", x"0976", x"08C4", x"07B3", x"0612", x"0412", x"01E6", x"FFC9", x"FE96", x"FE8A", x"FF2D", x"0060", x"0234", x"03F5", x"04CC", x"055A", x"0631", x"0703", x"07D2", x"08CD", x"0905", x"0802", x"0729", x"07B9", x"0983", x"0C6B", x"101F", x"1368", x"1510", x"155F", x"1464", x"11E1", x"0E6B", x"0B05", x"07F3", x"050F", x"02A9", x"0093", x"FE80", x"FCB3", x"FB94", x"FAE4", x"FA4A", x"F9CB", x"F954", x"F8FF", x"F918", x"FA01", x"FB45", x"FC2A", x"FC88", x"FC91", x"FC35", x"FBBE", x"FBC8", x"FC24", x"FC2F", x"FC42", x"FCA0", x"FC80", x"FB7C", x"FA83", x"F9FD", x"F95B", x"F924", x"F988", x"F911", x"F7D2", x"F7A1", x"F938", x"FBD4", x"FF98", x"040F", x"074B", x"08F2", x"09F0", x"0A06", x"0895", x"06C9", x"054F", x"03DF", x"0309", x"0352", x"0410", x"04AD", x"05D8", x"0761", x"08BA", x"09E9", x"0AE5", x"0B1C", x"0ACE", x"0AB4", x"0AD2", x"0AC0", x"0A27", x"08CF", x"0698", x"03C5", x"00ED", x"FEB9", x"FD0E", x"FBB7", x"FB0E", x"FAF8", x"FA77", x"F981", x"F910", x"F90C", x"F92D", x"F9F3", x"FAD4", x"FA5C", x"F933", x"F944", x"FABF", x"FD2C", x"00FE", x"050C", x"07BB", x"093C", x"0A3C", x"0A0D", x"08AD", x"0726", x"05AF", x"042A", x"0317", x"028B", x"0212", x"01B3", x"01E3", x"0272", x"030D", x"0354", x"0325", x"0281", x"01B9", x"0116", x"00E6", x"008A", x"FF5C", x"FD98", x"FB91", x"F906", x"F6B8", x"F570", x"F494", x"F3FB", x"F494", x"F5B8", x"F5EF", x"F5F1", x"F6B7", x"F79E", x"F8D2", x"FB20", x"FCB9", x"FC12", x"FADA", x"FA8A", x"FAD9", x"FC37", x"FF0C", x"0161", x"020E", x"0222", x"01B8", x"002D", x"FE2D", x"FCB3", x"FB7A", x"FAD8", x"FB83", x"FD26", x"FF2B", x"01AB", x"0496", x"075E", x"0989", x"0AEB", x"0B5A", x"0AFB", x"0A53", x"09DE", x"0988", x"08BB", x"072D", x"053E", x"02FC", x"00C5", x"FF7A", x"FF1F", x"FEEF", x"FF35", x"0047", x"0115", x"0130", x"0191", x"0243", x"02F9", x"0459", x"065B", x"0737", x"06B9", x"0675", x"071D", x"08B6", x"0BBB", x"0FA6", x"12B4", x"145E", x"152D", x"14D4", x"12FE", x"1050", x"0D63", x"0A34", x"0713", x"0457", x"01C5", x"FF17", x"FCA4", x"FAC4", x"F963", x"F822", x"F710", x"F61D", x"F551", x"F4E4", x"F553", x"F609", x"F663", x"F653", x"F61E", x"F592", x"F511", x"F55F", x"F5D4", x"F5FE", x"F69A", x"F7B1", x"F847", x"F871", x"F90A", x"F9B0", x"FA31", x"FB77", x"FCDD", x"FCA7", x"FB7E", x"FB2C", x"FBFC", x"FDF3", x"01C3", x"05FF", x"08A4", x"09D3", x"0A44", x"0957", x"0717", x"04D4", x"02C7", x"00CA", x"FFD8", x"0034", x"00E6", x"01B4", x"030E", x"0493", x"05CB", x"06E6", x"07A6", x"078F", x"0711", x"06CA", x"06BC", x"0663", x"0576", x"038D", x"0078", x"FC88", x"F89E", x"F53F", x"F247", x"EFCE", x"EE5D", x"ED80", x"EC5C", x"EB62", x"EAFD", x"EADC", x"EB59", x"ED29", x"EF05", x"EF8F", x"EFEB", x"F173", x"F3F7", x"F80E", x"FDC9", x"0325", x"0675", x"08A3", x"09F1", x"09D7", x"0909", x"0869", x"074C", x"05C9", x"04C4", x"03FC", x"02EF", x"0230", x"021B", x"0245", x"02BF", x"0355", x"03A9", x"038F", x"0384", x"03D0", x"0468", x"04E0", x"04A0", x"03B0", x"0222", x"002E", x"FEAE", x"FDE6", x"FD3A", x"FCB2", x"FD01", x"FD5A", x"FD1E", x"FD59", x"FE4B", x"FF3D", x"00EC", x"0383", x"04AE", x"0384", x"01D4", x"006F", x"FF69", x"003F", x"02C8", x"048E", x"0506", x"054F", x"04EA", x"036D", x"0208", x"00F5", x"FF78", x"FE6C", x"FE8F", x"FF47", x"004D", x"021A", x"0448", x"0643", x"07D3", x"08AF", x"086A", x"0753", x"0602", x"04EC", x"0405", x"02C4", x"00EA", x"FE9F", x"FBFD", x"F97C", x"F80F", x"F762", x"F6C8", x"F6C2", x"F76F", x"F7B4", x"F780", x"F7E3", x"F841", x"F89E", x"FA3D", x"FC8F", x"FD81", x"FD7C", x"FDF8", x"FF05", x"013D", x"05D2", x"0B3D", x"0F20", x"119E", x"131B", x"12BA", x"1107", x"0F07", x"0C67", x"08F0", x"059F", x"0296", x"FF2C", x"FBBE", x"F8BA", x"F623", x"F41C", x"F2F9", x"F241", x"F191", x"F0E5", x"F05C", x"F025", x"F035", x"F01F", x"EFEA", x"EF81", x"EEF5", x"EEB9", x"EF60", x"F03A", x"F0F9", x"F1FA", x"F2EB", x"F2DC", x"F26D", x"F21C", x"F162", x"F0C5", x"F14C", x"F1B2", x"F0A5", x"EF20", x"EE30", x"EDC2", x"EF1D", x"F2D3", x"F6D0", x"F975", x"FB57", x"FC4E", x"FBE9", x"FB32", x"FAE5", x"FA47", x"F97D", x"F986", x"F9F1", x"FA5F", x"FB55", x"FCC0", x"FE25", x"FF89", x"00EE", x"01B3", x"01E2", x"01DC", x"020A", x"027A", x"02F9", x"02EC", x"01E2", x"FFB8", x"FCA6", x"F978", x"F6D4", x"F453", x"F24B", x"F144", x"F09F", x"EFDF", x"EFC9", x"F04C", x"F0C2", x"F238", x"F4FC", x"F727", x"F7E9", x"F8B1", x"F9CC", x"FB87", x"FF9E", x"058C", x"0A6C", x"0D4D", x"0F06", x"0EF0", x"0D93", x"0CA4", x"0BFD", x"0A77", x"08E6", x"07D7", x"069B", x"0591", x"057B", x"05CB", x"0616", x"06D5", x"0781", x"0771", x"06E3", x"0633", x"056A", x"04D3", x"044B", x"0310", x"0107", x"FE39", x"FB0D", x"F883", x"F6E6", x"F5A2", x"F508", x"F541", x"F54A", x"F52B", x"F5B3", x"F65B", x"F6B8", x"F83C", x"FA42", x"FAA1", x"F980", x"F809", x"F5F1", x"F485", x"F5C7", x"F88E", x"FA9A", x"FC45", x"FD82", x"FD6C", x"FCFA", x"FD81", x"FDF0", x"FE05", x"FED2", x"0022", x"0160", x"0358", x"05FB", x"0866", x"0AAE", x"0CA3", x"0D7A", x"0D21", x"0C06", x"0A4A", x"0887", x"072E", x"05BC", x"041A", x"0281", x"0097", x"FEC1", x"FDD4", x"FD2F", x"FC4F", x"FC37", x"FCAF", x"FC97", x"FCC2", x"FD84", x"FDC4", x"FE35", x"0062", x"02CB", x"03B6", x"0430", x"0451", x"03C7", x"04BE", x"085B", x"0C39", x"0EED", x"10E4", x"1123", x"0F77", x"0DAD", x"0C40", x"09F8", x"074D", x"04C5", x"018A", x"FDE9", x"FAC0", x"F7E0", x"F52D", x"F364", x"F25A", x"F16F", x"F0D7", x"F050", x"EFCA", x"EFB6", x"F01A", x"F07F", x"F0CA", x"F0CC", x"F035", x"EFC6", x"F028", x"F085", x"F137", x"F296", x"F3A3", x"F3EB", x"F43F", x"F42C", x"F2FB", x"F227", x"F24D", x"F1CD", x"F096", x"EFB3", x"EEAD", x"EE31", x"F079", x"F52F", x"F9ED", x"FE16", x"012E", x"01F9", x"015D", x"0130", x"0131", x"00D2", x"00AC", x"0068", x"FF59", x"FE77", x"FE48", x"FE5D", x"FEC3", x"FFA3", x"004D", x"006A", x"0064", x"002E", x"0004", x"0044", x"00A0", x"0069", x"FF66", x"FD35", x"FA06", x"F700", x"F454", x"F1C7", x"EFEF", x"EEDE", x"EDA0", x"EC97", x"EC57", x"EBD5", x"EB24", x"EBBA", x"ED4F", x"EE60", x"EF8A", x"F109", x"F21D", x"F41D", x"F8BB", x"FE8E", x"037F", x"076E", x"09A2", x"0949", x"085A", x"082D", x"07F8", x"0761", x"071C", x"0663", x"051E", x"0469", x"0493", x"04BC", x"0565", x"068D", x"077F", x"080B", x"0883", x"08AA", x"08AA", x"08F3", x"0937", x"08ED", x"07E7", x"05CB", x"0335", x"0108", x"FF48", x"FDD9", x"FD60", x"FD71", x"FD69", x"FE0A", x"FF5A", x"0006", x"008A", x"020A", x"032A", x"02F6", x"0244", x"00BC", x"FE07", x"FC83", x"FDAC", x"FFC8", x"01EA", x"0409", x"04C1", x"0393", x"02A1", x"0257", x"01C8", x"0180", x"01EC", x"01FE", x"0222", x"033B", x"04D0", x"0647", x"0830", x"09EB", x"0AB1", x"0AA4", x"09D5", x"082B", x"0658", x"04F6", x"03B3", x"02A1", x"0189", x"0008", x"FEE4", x"FE81", x"FE6F", x"FEC7", x"0004", x"0123", x"01B6", x"02AC", x"034E", x"02E4", x"0306", x"0477", x"059F", x"064A", x"06EE", x"0671", x"052E", x"0601", x"0917", x"0C99", x"1038", x"1324", x"13B7", x"12A3", x"1205", x"1183", x"10B5", x"1024", x"0F07", x"0C64", x"0931", x"0627", x"0304", x"006E", x"FEEC", x"FDC3", x"FC8D", x"FB95", x"FA49", x"F8DB", x"F7FA", x"F793", x"F774", x"F79E", x"F791", x"F71A", x"F72D", x"F7C5", x"F870", x"F9B3", x"FB6B", x"FC5C", x"FCCA", x"FD52", x"FCB5", x"FB0C", x"FA21", x"F9C3", x"F8BF", x"F7D8", x"F715", x"F562", x"F448", x"F601", x"F994", x"FD9B", x"01DF", x"04E1", x"0565", x"04F0", x"04FF", x"04FA", x"052B", x"05E8", x"062A", x"058B", x"0510", x"04D9", x"046D", x"0468", x"04B4", x"04BE", x"0495", x"04B3", x"04D4", x"055C", x"0671", x"07BA", x"08A7", x"08C5", x"078B", x"0577", x"035A", x"012D", x"FF31", x"FDE5", x"FCBB", x"FB3C", x"FA5A", x"F9FD", x"F90E", x"F84C", x"F8B9", x"F971", x"FA19", x"FB81", x"FCC8", x"FD3B", x"FEA4", x"0203", x"05F4", x"09D4", x"0D5E", x"0ED5", x"0DF2", x"0CA8", x"0B8C", x"0A59", x"09A0", x"094B", x"0824", x"068C", x"0545", x"0428", x"033C", x"0328", x"0364", x"0373", x"0396", x"03A3", x"0349", x"02E7", x"02A3", x"01FE", x"00FE", x"FF5B", x"FCB0", x"F9A9", x"F707", x"F4A1", x"F2F6", x"F2A9", x"F2DC", x"F336", x"F46D", x"F5E1", x"F684", x"F794", x"F9BE", x"FB7F", x"FC8A", x"FD41", x"FC50", x"F9D9", x"F8A6", x"F9B3", x"FBC5", x"FEB6", x"01DC", x"0309", x"023F", x"0162", x"0083", x"FFA3", x"FFBE", x"00B7", x"017F", x"0297", x"0468", x"0643", x"0839", x"0AA8", x"0CC4", x"0E0D", x"0EB5", x"0E6F", x"0D69", x"0C6B", x"0BC0", x"0B4A", x"0AF0", x"0A07", x"0845", x"066B", x"04C8", x"0344", x"02AA", x"02E6", x"02DC", x"02E0", x"037F", x"039B", x"0331", x"03EF", x"05AC", x"072C", x"08FD", x"0A87", x"0A10", x"08C9", x"0910", x"0AB2", x"0D24", x"1084", x"131E", x"133D", x"120C", x"10D1", x"0F4A", x"0E21", x"0DA9", x"0C6A", x"09FB", x"0736", x"0423", x"00F2", x"FEC3", x"FD4A", x"FBCB", x"FA91", x"F9A0", x"F863", x"F780", x"F759", x"F739", x"F71D", x"F752", x"F710", x"F69C", x"F72B", x"F84E", x"F9BF", x"FC32", x"FF00", x"00CE", x"0251", x"0396", x"0329", x"01C5", x"0125", x"0098", x"FF9B", x"FF10", x"FE3F", x"FBE5", x"FA41", x"FB10", x"FD81", x"0132", x"05F1", x"099E", x"0B12", x"0B8F", x"0BAA", x"0B12", x"0AC6", x"0B08", x"0B00", x"0AB0", x"0A7B", x"09FB", x"0938", x"08D1", x"0866", x"07E6", x"0784", x"0727", x"06C2", x"06E9", x"076D", x"07D6", x"0802", x"073C", x"04DF", x"01CE", x"FEB0", x"FB5C", x"F88C", x"F6DA", x"F528", x"F37D", x"F2C4", x"F215", x"F0A0", x"EFA5", x"EFD8", x"F04A", x"F1A3", x"F43E", x"F63C", x"F74B", x"F952", x"FCAB", x"009F", x"05A7", x"0AB0", x"0D9E", x"0E7F", x"0E78", x"0DB0", x"0CE4", x"0D29", x"0DF1", x"0E4C", x"0E83", x"0E35", x"0D04", x"0BE2", x"0B1C", x"0A1F", x"0952", x"08FC", x"0875", x"0802", x"084D", x"08AE", x"08C3", x"0901", x"08B2", x"0751", x"05DA", x"04A7", x"0348", x"02AD", x"034B", x"03D8", x"0436", x"04F7", x"04E3", x"03A8", x"0328", x"03AB", x"0425", x"04DE", x"0558", x"03D1", x"00EB", x"FF33", x"FF2F", x"0073", x"0358", x"0665", x"0797", x"0730", x"061F", x"0478", x"0302", x"02B3", x"032A", x"03EB", x"0504", x"0621", x"06F7", x"081D", x"0943", x"0A08", x"0A61", x"09FD", x"08B9", x"074F", x"0643", x"055B", x"04BE", x"0449", x"02F6", x"00F3", x"FF24", x"FD4D", x"FBAD", x"FB33", x"FB4F", x"FB24", x"FB9E", x"FCA0", x"FD06", x"FD6B", x"FF21", x"013F", x"038D", x"0688", x"08BD", x"08A2", x"07E5", x"080F", x"0907", x"0B66", x"0F26", x"1214", x"12F7", x"12A6", x"1162", x"0F66", x"0DFD", x"0D38", x"0C1E", x"0AA0", x"08C1", x"05F3", x"02D8", x"0030", x"FD82", x"FACB", x"F896", x"F66E", x"F45F", x"F335", x"F2BD", x"F243", x"F217", x"F20B", x"F15E", x"F0BF", x"F0E3", x"F145", x"F206", x"F3D3", x"F585", x"F689", x"F788", x"F7F0", x"F6B1", x"F50B", x"F40B", x"F31E", x"F2B3", x"F344", x"F318", x"F16A", x"F000", x"EFF0", x"F10D", x"F400", x"F864", x"FC1A", x"FE45", x"FF7E", x"FFC3", x"FF61", x"FF7D", x"008A", x"0206", x"03C8", x"0548", x"05F4", x"05E7", x"0570", x"04CF", x"0451", x"0405", x"03A2", x"0360", x"037C", x"0393", x"03B4", x"03CE", x"031F", x"016E", x"FF7C", x"FD61", x"FB1F", x"F99D", x"F8DA", x"F7E2", x"F72A", x"F71A", x"F6B9", x"F5DA", x"F5CA", x"F681", x"F79A", x"F9E2", x"FCD9", x"FE77", x"FED8", x"FF8F", x"00F2", x"0349", x"0744", x"0BB3", x"0E87", x"0FA6", x"0F91", x"0E46", x"0CA1", x"0BDA", x"0BC6", x"0BFF", x"0C6B", x"0C67", x"0B90", x"0A54", x"0900", x"0784", x"065C", x"0571", x"0482", x"03E7", x"03D4", x"03C0", x"0386", x"031A", x"01C4", x"FF5D", x"FCD4", x"FA5E", x"F849", x"F77F", x"F7DE", x"F872", x"F92E", x"FA36", x"FA4C", x"F9C6", x"F9D8", x"FA5C", x"FADC", x"FBD0", x"FC4A", x"FAB1", x"F813", x"F67B", x"F64E", x"F7F3", x"FBB2", x"FFCD", x"023C", x"034E", x"037F", x"02CF", x"0210", x"0283", x"03BB", x"0574", x"079F", x"099E", x"0AE0", x"0B9F", x"0BEF", x"0BAF", x"0B13", x"0A16", x"08A2", x"0731", x"05E8", x"04AC", x"03AC", x"02C6", x"016E", x"FFD7", x"FE75", x"FD24", x"FC43", x"FC4D", x"FC95", x"FCA3", x"FCFF", x"FD66", x"FD22", x"FD1D", x"FE12", x"FF3E", x"0105", x"0393", x"0536", x"04A3", x"0369", x"0279", x"0216", x"0361", x"0683", x"0916", x"0A23", x"0A35", x"0914", x"06A2", x"0469", x"02C1", x"0142", x"0027", x"FF8B", x"FE6D", x"FCCF", x"FAF4", x"F8C5", x"F667", x"F46F", x"F2BD", x"F147", x"F099", x"F06D", x"F070", x"F0E2", x"F168", x"F17C", x"F199", x"F1FB", x"F257", x"F33C", x"F4EF", x"F66D", x"F795", x"F8CC", x"F920", x"F804", x"F6BC", x"F593", x"F426", x"F3A7", x"F420", x"F37B", x"F174", x"EFDE", x"EF37", x"EFEC", x"F363", x"F893", x"FCC0", x"FF5B", x"00E6", x"00CF", x"FF95", x"FEE9", x"FEEE", x"FF4A", x"0051", x"01A8", x"021B", x"018E", x"005E", x"FEB3", x"FD02", x"FBB6", x"FAA4", x"F9DA", x"F95B", x"F8FB", x"F8AD", x"F87A", x"F7A2", x"F612", x"F430", x"F1F6", x"EF9D", x"EE2E", x"ED4D", x"EC39", x"EB6E", x"EAE5", x"E9A8", x"E832", x"E7D4", x"E82C", x"E956", x"EC69", x"F010", x"F20F", x"F2D0", x"F380", x"F421", x"F5D7", x"F9D2", x"FE52", x"0151", x"0337", x"043C", x"03F2", x"038D", x"042D", x"0583", x"0746", x"09CD", x"0C22", x"0D81", x"0DDB", x"0D74", x"0C4E", x"0AF8", x"097E", x"07FB", x"06C5", x"05F1", x"0535", x"04CF", x"0458", x"031A", x"0172", x"FFD9", x"FE0B", x"FC91", x"FC24", x"FC06", x"FBAB", x"FBD8", x"FBFE", x"FB23", x"FA23", x"F9BA", x"F91B", x"F8F3", x"FA16", x"FAA5", x"F920", x"F6E5", x"F4F6", x"F37D", x"F44A", x"F7C6", x"FB4F", x"FD49", x"FE5C", x"FE1B", x"FC64", x"FAD2", x"FA63", x"FA8F", x"FBD4", x"FE8D", x"0185", x"03C3", x"052E", x"0598", x"04FC", x"03E7", x"02A8", x"0141", x"0016", x"FF0B", x"FE33", x"FDB4", x"FD23", x"FC3F", x"FB69", x"FAC5", x"FA12", x"FA0F", x"FAD3", x"FB87", x"FC3A", x"FD9A", x"FEA5", x"FF19", x"FFF0", x"00FB", x"0195", x"0322", x"05B1", x"0703", x"068C", x"059C", x"041A", x"030A", x"04B2", x"089E", x"0C3B", x"0F00", x"1110", x"115E", x"1058", x"0F91", x"0EF9", x"0E18", x"0DB8", x"0D9E", x"0C9F", x"0A8D", x"077F", x"038D", x"FF35", x"FB18", x"F75B", x"F452", x"F23A", x"F0C3", x"F040", x"F06A", x"F075", x"F047", x"F080", x"F0AC", x"F0E9", x"F22F", x"F3BF", x"F4A9", x"F592", x"F691", x"F635", x"F515", x"F43B", x"F2DA", x"F15F", x"F1BD", x"F2F3", x"F2AA", x"F16F", x"EFFD", x"EE26", x"EDEA", x"F181", x"F6DE", x"FB81", x"FF4B", x"0193", x"0155", x"001A", x"FF5F", x"FEB8", x"FE6F", x"FF7B", x"012B", x"026C", x"0306", x"030D", x"0256", x"0188", x"00DC", x"0066", x"0023", x"FFF8", x"0009", x"00A4", x"013D", x"012C", x"00B5", x"FFDF", x"FE3D", x"FCC8", x"FBF5", x"FAE2", x"F97B", x"F8C3", x"F814", x"F6DB", x"F630", x"F601", x"F547", x"F55A", x"F73C", x"F934", x"FA0A", x"FA7C", x"F9F2", x"F8D0", x"F98C", x"FD27", x"016C", x"054E", x"087A", x"09CA", x"0913", x"07F4", x"06F8", x"05FF", x"05C2", x"0674", x"075D", x"07AA", x"071B", x"0586", x"0365", x"0115", x"FED3", x"FD22", x"FC20", x"FB55", x"FB1A", x"FB2D", x"FA78", x"F893", x"F67E", x"F423", x"F1BD", x"F08E", x"F071", x"F012", x"EFE2", x"F05B", x"F073", x"F021", x"F08F", x"F0E8", x"F0D0", x"F1CF", x"F41E", x"F5AD", x"F627", x"F600", x"F48E", x"F2DF", x"F385", x"F66A", x"F987", x"FC55", x"FE87", x"FEFD", x"FE26", x"FDA5", x"FDA6", x"FE34", x"001D", x"039C", x"076E", x"0AAD", x"0CF4", x"0E09", x"0DFC", x"0D1B", x"0BCE", x"0A2C", x"0832", x"0646", x"052A", x"0485", x"03AA", x"02B1", x"01A6", x"0029", x"FEFD", x"FEF4", x"FF61", x"FFAB", x"0066", x"014B", x"0195", x"0200", x"0307", x"038D", x"03F3", x"0583", x"074E", x"07E6", x"0788", x"060B", x"0322", x"00DC", x"016C", x"03F5", x"06D2", x"09AB", x"0B3F", x"0A83", x"08A0", x"06DD", x"0530", x"0404", x"0431", x"0519", x"0593", x"04F6", x"0311", x"FFDD", x"FC0D", x"F83A", x"F4E2", x"F226", x"F002", x"EEBC", x"EEBF", x"EF77", x"F030", x"F115", x"F221", x"F2ED", x"F467", x"F71D", x"FA1A", x"FCE6", x"FFF4", x"0247", x"02FC", x"02F8", x"0269", x"00A3", x"FEFC", x"FEE3", x"FF28", x"FEBB", x"FE20", x"FCBC", x"FA5A", x"F98E", x"FBC9", x"FF5A", x"0320", x"06E3", x"090A", x"08FE", x"0848", x"07B4", x"06D6", x"0699", x"07D6", x"09B8", x"0B27", x"0BD4", x"0B58", x"0997", x"0754", x"0537", x"0364", x"01BC", x"002B", x"FF2A", x"FECB", x"FE87", x"FE13", x"FD92", x"FC6F", x"FAAD", x"F947", x"F834", x"F6AD", x"F51E", x"F3FD", x"F26D", x"F0CC", x"F03D", x"F00B", x"EFDE", x"F123", x"F3EB", x"F688", x"F8B4", x"FA71", x"FA60", x"F974", x"FA87", x"FDE6", x"0246", x"0755", x"0C1D", x"0E98", x"0F37", x"0F61", x"0F0D", x"0E43", x"0E5F", x"0F9B", x"10FB", x"1261", x"133F", x"12DC", x"115A", x"0F83", x"0D9C", x"0C13", x"0B1D", x"0A90", x"0A90", x"0AE0", x"0ACC", x"0A09", x"08D6", x"06F9", x"04E2", x"0393", x"02F5", x"0296", x"02AA", x"030D", x"02A5", x"01CD", x"0115", x"FFED", x"FEB2", x"FED6", x"FFF8", x"00DF", x"018B", x"017B", x"FFB8", x"FDD3", x"FE13", x"001D", x"02FA", x"0661", x"08EB", x"0922", x"081A", x"0714", x"05FE", x"056B", x"0686", x"08FA", x"0BA5", x"0E46", x"1011", x"106B", x"0F98", x"0E71", x"0D0D", x"0B9E", x"0A18", x"0898", x"0750", x"062A", x"04F0", x"039C", x"0219", x"0043", x"FEA3", x"FE03", x"FDEE", x"FE75", x"FFD9", x"0197", x"02FF", x"04C1", x"06C0", x"081C", x"09AA", x"0C44", x"0EE2", x"10B6", x"11E4", x"1143", x"0E3E", x"0B80", x"0AE9", x"0BE1", x"0E31", x"11A0", x"13D1", x"13CC", x"1313", x"121C", x"1032", x"0E94", x"0E29", x"0DE5", x"0D72", x"0D03", x"0B6D", x"07FC", x"03D1", x"FF9C", x"FB6E", x"F812", x"F5C7", x"F427", x"F326", x"F2DB", x"F2AB", x"F271", x"F24D", x"F1F7", x"F1D8", x"F271", x"F37A", x"F4C3", x"F673", x"F7AE", x"F7FF", x"F7F0", x"F765", x"F60D", x"F52E", x"F578", x"F5D5", x"F610", x"F641", x"F524", x"F304", x"F284", x"F477", x"F7AF", x"FC27", x"00E5", x"038D", x"0432", x"0494", x"0485", x"03E7", x"0451", x"05E8", x"07B1", x"09D4", x"0C14", x"0CFA", x"0C4A", x"0ACE", x"0891", x"05F1", x"03B1", x"0200", x"00D8", x"00B4", x"0107", x"015B", x"01B4", x"019A", x"00E2", x"0062", x"0044", x"FFDB", x"FFDD", x"0053", x"0029", x"FF9C", x"FF71", x"FEAD", x"FD78", x"FDAA", x"FF3A", x"00A3", x"026E", x"03AF", x"0272", x"0043", x"0011", x"01DB", x"051E", x"0A63", x"0F6E", x"11C4", x"12A0", x"1316", x"125D", x"112F", x"112D", x"1169", x"1167", x"120E", x"1275", x"1165", x"0F5D", x"0D0B", x"0A10", x"076D", x"05AD", x"045E", x"036F", x"0316", x"0289", x"01B9", x"00FC", x"FFF4", x"FEAF", x"FE09", x"FD93", x"FD14", x"FD25", x"FD83", x"FD35", x"FCED", x"FCCB", x"FBE0", x"FB04", x"FBB5", x"FD16", x"FEAB", x"00D5", x"01ED", x"00C3", x"FF82", x"FFCD", x"0148", x"045C", x"08D7", x"0C05", x"0CC5", x"0C94", x"0BC1", x"0A45", x"09EC", x"0B3B", x"0D2C", x"0FD9", x"132E", x"158A", x"165D", x"15E6", x"13F8", x"10BD", x"0D82", x"0A6F", x"07BC", x"0619", x"0529", x"042A", x"037D", x"02E6", x"01CF", x"0112", x"013A", x"014E", x"01A6", x"02E4", x"03EF", x"048D", x"05D6", x"06F9", x"06EB", x"0731", x"0851", x"08EF", x"0991", x"0A6D", x"0920", x"05B4", x"02FE", x"01B8", x"0190", x"03A8", x"06E5", x"0815", x"079E", x"0708", x"05C2", x"0415", x"03A6", x"03BB", x"032B", x"0322", x"0379", x"02C9", x"013E", x"FF5A", x"FC7B", x"F932", x"F6C2", x"F4E9", x"F3A1", x"F356", x"F36B", x"F33A", x"F32A", x"F2D7", x"F224", x"F217", x"F307", x"F45C", x"F6B3", x"F9C6", x"FC0B", x"FDC1", x"FF49", x"FF81", x"FE80", x"FE33", x"FE45", x"FE2B", x"FEDF", x"FF70", x"FD78", x"FA62", x"F864", x"F799", x"F8A6", x"FCA1", x"00D5", x"02DC", x"03C8", x"0414", x"032F", x"02B8", x"03BC", x"04C0", x"05BE", x"078F", x"08FF", x"0941", x"08F3", x"078A", x"046E", x"00EE", x"FD81", x"F9FE", x"F786", x"F65E", x"F569", x"F4D5", x"F4BA", x"F3CB", x"F266", x"F1B3", x"F0BF", x"EF53", x"EED8", x"EEA5", x"EDDB", x"EE08", x"EF1B", x"EF05", x"EED5", x"F016", x"F17F", x"F336", x"F685", x"F8C9", x"F7FA", x"F68D", x"F5F3", x"F609", x"F8CB", x"FE8F", x"03BE", x"06F5", x"09A5", x"0B04", x"0B1E", x"0C2A", x"0E15", x"0F54", x"10C0", x"12A1", x"1346", x"12F3", x"1250", x"1051", x"0D56", x"0AE3", x"08C2", x"06F5", x"069E", x"06BC", x"0610", x"053C", x"03DE", x"0147", x"FF03", x"FE01", x"FCEB", x"FC4A", x"FCCC", x"FCC5", x"FC26", x"FC7B", x"FC8B", x"FB1C", x"FA16", x"F9C5", x"F90F", x"F967", x"FB2C", x"FB56", x"F9BC", x"F876", x"F77D", x"F732", x"F9B2", x"FD92", x"FFE0", x"00FC", x"0159", x"0024", x"FEE8", x"FF5E", x"004C", x"014E", x"0361", x"0548", x"0664", x"07BB", x"08B1", x"0808", x"06BE", x"0506", x"022E", x"FFC5", x"FEE1", x"FE1D", x"FD91", x"FDE3", x"FD93", x"FC8E", x"FCD2", x"FDC8", x"FE47", x"FF99", x"0175", x"020B", x"02C7", x"04C1", x"05E8", x"0633", x"07A3", x"0917", x"0A09", x"0C68", x"0EF3", x"0EAC", x"0CD7", x"0B1B", x"090D", x"086F", x"0B08", x"0E41", x"0FEE", x"10F4", x"10D1", x"0EF6", x"0D92", x"0D5B", x"0CC6", x"0C28", x"0C0F", x"0B0B", x"0938", x"07A1", x"0548", x"01BD", x"FE3B", x"FA8E", x"F696", x"F3F6", x"F2D6", x"F1F5", x"F1C9", x"F235", x"F1A6", x"F0E4", x"F11E", x"F144", x"F148", x"F25D", x"F356", x"F340", x"F3BC", x"F475", x"F386", x"F229", x"F17B", x"F05E", x"EFE2", x"F198", x"F350", x"F32C", x"F2E3", x"F29D", x"F242", x"F3EF", x"F839", x"FC0E", x"FEC2", x"00D8", x"0142", x"0068", x"0078", x"011F", x"0180", x"02A5", x"043D", x"0527", x"0630", x"0792", x"07BC", x"06E5", x"05B5", x"034B", x"0067", x"FECC", x"FDD5", x"FCC8", x"FC96", x"FC3F", x"FABE", x"F9AD", x"F9CB", x"F986", x"F9AC", x"FAB1", x"FAA2", x"F98E", x"F982", x"F942", x"F7DC", x"F739", x"F769", x"F708", x"F7D3", x"FA3D", x"FB31", x"FA14", x"F8F7", x"F787", x"F6A1", x"F91F", x"FE11", x"025D", x"0601", x"08BD", x"0930", x"08BC", x"0944", x"09A0", x"0963", x"09D3", x"09BF", x"08A6", x"0802", x"0772", x"0575", x"02EF", x"002C", x"FC4D", x"F8C3", x"F711", x"F5DA", x"F4C9", x"F4A2", x"F3DF", x"F1F0", x"F09E", x"EFCA", x"EE60", x"EDD9", x"EE3D", x"EDE6", x"EDC7", x"EED5", x"EF48", x"EF01", x"EFA6", x"F05B", x"F0AF", x"F293", x"F526", x"F5DC", x"F56B", x"F4E2", x"F3AA", x"F392", x"F68E", x"FA82", x"FDC3", x"00AE", x"023E", x"01EC", x"022D", x"039B", x"051D", x"0734", x"09D0", x"0AF1", x"0B0C", x"0B59", x"0A92", x"088A", x"066E", x"0387", x"FF5E", x"FC50", x"FA9B", x"F8FA", x"F850", x"F8B9", x"F856", x"F7D4", x"F8B8", x"F9A4", x"FA70", x"FC7E", x"FE89", x"FF72", x"0116", x"033C", x"0401", x"046F", x"0548", x"04CE", x"03FF", x"04C0", x"04FF", x"031A", x"00A8", x"FD9E", x"F9CD", x"F847", x"FA06", x"FC6D", x"FED7", x"0158", x"0224", x"0155", x"013C", x"013B", x"0086", x"0036", x"FFF9", x"FE7E", x"FD38", x"FCBC", x"FB6C", x"F97E", x"F7B8", x"F4E7", x"F1B0", x"F01E", x"EFAE", x"EF99", x"F0A3", x"F215", x"F264", x"F2E7", x"F40E", x"F4C5", x"F5B8", x"F7B7", x"F930", x"F9FE", x"FBBB", x"FD15", x"FD3D", x"FD95", x"FDF3", x"FD21", x"FCF7", x"FE0D", x"FE00", x"FC6B", x"FAAB", x"F821", x"F5BF", x"F636", x"F91A", x"FC30", x"FF77", x"0254", x"035C", x"03B8", x"04CA", x"05BC", x"06AC", x"0838", x"0923", x"08FA", x"0915", x"08EF", x"07B8", x"063B", x"0422", x"004C", x"FC79", x"F9FD", x"F7FA", x"F6C2", x"F6D5", x"F648", x"F489", x"F355", x"F252", x"F0EA", x"F0AC", x"F165", x"F131", x"F121", x"F21D", x"F24A", x"F1D0", x"F24D", x"F291", x"F264", x"F423", x"F719", x"F88C", x"F8F2", x"F8D7", x"F768", x"F69A", x"F931", x"FD86", x"01D5", x"065B", x"098B", x"0A61", x"0AE0", x"0C0F", x"0CF5", x"0E64", x"1086", x"1196", x"11C9", x"126A", x"126C", x"115F", x"106A", x"0E9C", x"0B4B", x"0870", x"0697", x"046E", x"0295", x"0171", x"FF59", x"FCBD", x"FB2D", x"F9CF", x"F84B", x"F818", x"F873", x"F854", x"F8F2", x"FA3A", x"FA7A", x"FA7B", x"FAE4", x"FA6E", x"F9C9", x"FAB9", x"FB94", x"FB29", x"FA61", x"F8D6", x"F640", x"F533", x"F6DD", x"F96C", x"FC8C", x"FFE6", x"0175", x"0158", x"0185", x"01DD", x"0220", x"0392", x"0525", x"0558", x"0595", x"0636", x"05FB", x"0580", x"053F", x"0374", x"008B", x"FEBB", x"FD6D", x"FBEA", x"FB88", x"FB76", x"FA5A", x"F9B8", x"FA46", x"FAC5", x"FBF4", x"FE92", x"00F4", x"02DE", x"05C3", x"0852", x"09CD", x"0B9E", x"0D41", x"0D38", x"0D96", x"0EFD", x"0F4D", x"0E65", x"0D41", x"0A5C", x"067B", x"0503", x"05C9", x"06FA", x"08E8", x"0A90", x"09D0", x"0815", x"0744", x"0669", x"059C", x"05CF", x"0578", x"03DB", x"02C1", x"01F6", x"004B", x"FEA9", x"FCDE", x"F99A", x"F60C", x"F3CC", x"F203", x"F0C9", x"F0EE", x"F130", x"F0C3", x"F0CF", x"F0F6", x"F093", x"F0EE", x"F1FD", x"F273", x"F2E5", x"F3C6", x"F389", x"F2C8", x"F2A7", x"F1F7", x"F0A8", x"F0EC", x"F22B", x"F29B", x"F2DA", x"F298", x"F061", x"EE3A", x"EEE6", x"F184", x"F525", x"FA0E", x"FE42", x"0051", x"01E7", x"03B5", x"04DE", x"0627", x"07CB", x"0833", x"07CE", x"07BC", x"0767", x"06AF", x"068C", x"05EE", x"03FB", x"024A", x"0112", x"FF8E", x"FEB0", x"FE83", x"FD70", x"FBC1", x"FACB", x"F999", x"F878", x"F8C0", x"F966", x"F949", x"F9CC", x"FAA5", x"FA85", x"FA9B", x"FB79", x"FB5F", x"FB1C", x"FC9D", x"FE56", x"FED4", x"FF1D", x"FE58", x"FBBD", x"FA5F", x"FC3D", x"FFB4", x"041B", x"0951", x"0CEA", x"0E4B", x"0F6D", x"1084", x"10D7", x"11AC", x"12AB", x"1286", x"11E9", x"118C", x"1057", x"0ECD", x"0D8E", x"0B80", x"0878", x"0634", x"0465", x"0272", x"016C", x"00D8", x"FF1E", x"FD38", x"FBD6", x"F9F3", x"F82D", x"F795", x"F718", x"F65E", x"F6CD", x"F780", x"F78A", x"F830", x"F942", x"F97E", x"FA73", x"FD0A", x"FF51", x"00B9", x"01D7", x"0132", x"FF05", x"FE8B", x"0057", x"030D", x"06DB", x"0AF5", x"0D05", x"0DCD", x"0F02", x"1002", x"10DF", x"1279", x"136D", x"12AE", x"11C0", x"109F", x"0EC2", x"0D70", x"0CAB", x"0AAB", x"0830", x"0683", x"0489", x"0286", x"01C0", x"010C", x"FFAF", x"FF57", x"000F", x"0087", x"01DF", x"0439", x"05F4", x"07BB", x"0A84", x"0CCB", x"0E39", x"1001", x"10C7", x"0FEC", x"0F9C", x"0FBA", x"0E64", x"0C33", x"094A", x"03E8", x"FE07", x"FAFC", x"FA6B", x"FB5C", x"FE52", x"0129", x"01A9", x"016A", x"0173", x"00B2", x"0008", x"0031", x"FFA2", x"FE50", x"FDD2", x"FD7A", x"FCE8", x"FD34", x"FD8F", x"FC96", x"FB87", x"FAEF", x"F9DD", x"F941", x"F9C5", x"F9E5", x"F9B0", x"FA53", x"FAF1", x"FB35", x"FC61", x"FDDB", x"FEAA", x"FFFE", x"01D1", x"02AE", x"0380", x"048A", x"040D", x"029B", x"0211", x"0168", x"FFE8", x"FED3", x"FD02", x"F926", x"F60D", x"F5C9", x"F71D", x"FA2E", x"FEF8", x"02C7", x"048D", x"0665", x"0843", x"093E", x"0A88", x"0BC8", x"0B88", x"0A71", x"099F", x"0822", x"0663", x"0538", x"036D", x"0091", x"FDFE", x"FB5A", x"F84E", x"F601", x"F44B", x"F1EC", x"EFEA", x"EEC5", x"EDAD", x"ED14", x"EDEC", x"EEC7", x"EF7C", x"F10A", x"F298", x"F35F", x"F4DC", x"F689", x"F70B", x"F7DC", x"F9EA", x"FB5D", x"FC60", x"FD94", x"FD11", x"FAB7", x"F9F1", x"FBA2", x"FEA8", x"03A4", x"09A3", x"0D98", x"0FCA", x"1208", x"13B6", x"14B1", x"164A", x"1796", x"1786", x"1748", x"1728", x"164A", x"159D", x"1563", x"1441", x"1269", x"10B4", x"0E4C", x"0B6F", x"0954", x"0738", x"0486", x"0281", x"00F6", x"FF0A", x"FDD4", x"FD89", x"FCF3", x"FCC3", x"FDBC", x"FE94", x"FF25", x"007A", x"0131", x"0091", x"0096", x"0130", x"0108", x"00D8", x"0080", x"FDD3", x"FA10", x"F83C", x"F83E", x"F9A3", x"FD1C", x"00B4", x"0232", x"02CF", x"03D9", x"047B", x"0565", x"071B", x"0819", x"07E8", x"0790", x"06BD", x"0571", x"04FC", x"04ED", x"044B", x"03D4", x"0353", x"020C", x"0103", x"00C9", x"0012", x"FF40", x"FF55", x"FF6D", x"FF8A", x"00F4", x"02DC", x"0423", x"0627", x"08C4", x"0ABC", x"0D18", x"102C", x"1216", x"1315", x"14D4", x"1636", x"1674", x"16B8", x"15AA", x"11AE", x"0D40", x"0A76", x"08D8", x"08C3", x"0AAF", x"0BF9", x"0B8E", x"0B3D", x"0B1C", x"0ABA", x"0B03", x"0BD9", x"0BAD", x"0AF7", x"0A2B", x"08C1", x"0742", x"0695", x"0599", x"040C", x"0286", x"006D", x"FDA0", x"FBC2", x"FA77", x"F8D0", x"F789", x"F6EA", x"F5C7", x"F4DF", x"F511", x"F4E3", x"F43F", x"F451", x"F473", x"F40D", x"F48A", x"F55A", x"F50F", x"F4CE", x"F590", x"F610", x"F69B", x"F7B8", x"F778", x"F533", x"F376", x"F325", x"F3FE", x"F6ED", x"FB7A", x"FF22", x"01C5", x"0481", x"06C0", x"08A6", x"0AEC", x"0CFB", x"0DDB", x"0E33", x"0DD7", x"0C87", x"0B5E", x"0AB0", x"09B2", x"08C5", x"07E2", x"061D", x"03E8", x"0256", x"0075", x"FE2C", x"FC61", x"FAC2", x"F8B8", x"F78B", x"F74D", x"F6C4", x"F6B7", x"F7C4", x"F8C6", x"F9F7", x"FC2C", x"FE02", x"FEB0", x"FFC0", x"0114", x"01B1", x"0289", x"0350", x"01D9", x"FEDF", x"FCE9", x"FC1C", x"FCDE", x"0030", x"047E", x"073F", x"0942", x"0B0C", x"0BF5", x"0C91", x"0DA9", x"0DDB", x"0CCF", x"0B81", x"09B8", x"0772", x"05EC", x"050A", x"03ED", x"030D", x"0251", x"00D1", x"FF22", x"FDEC", x"FC2C", x"F9FF", x"F850", x"F68A", x"F492", x"F390", x"F338", x"F2B9", x"F2EB", x"F3C3", x"F418", x"F481", x"F570", x"F5A9", x"F576", x"F659", x"F79C", x"F8C3", x"FAAE", x"FC1F", x"FB49", x"F9C3", x"F939", x"F989", x"FB7A", x"FFA8", x"03C9", x"0647", x"085F", x"0A24", x"0B0D", x"0C2C", x"0D73", x"0D64", x"0C39", x"0A9A", x"083D", x"05C7", x"0459", x"0373", x"0297", x"024E", x"01BA", x"0079", x"FF78", x"FEBD", x"FD5B", x"FC36", x"FBB2", x"FAED", x"FAB9", x"FBED", x"FD57", x"FEB3", x"0102", x"035D", x"0530", x"07A9", x"0A46", x"0B3A", x"0B7A", x"0BD7", x"0B28", x"09DE", x"0932", x"06FF", x"0271", x"FDE7", x"FA83", x"F818", x"F846", x"FAF1", x"FD36", x"FE68", x"FFB1", x"005D", x"004B", x"00C4", x"0149", x"00AF", x"FFD3", x"FEE7", x"FD6D", x"FC49", x"FC1B", x"FC46", x"FCD8", x"FE10", x"FEC9", x"FECB", x"FEE2", x"FE62", x"FD1C", x"FC27", x"FB4C", x"FA19", x"F975", x"F99A", x"F966", x"F967", x"FA3D", x"FAF4", x"FB7A", x"FCDF", x"FDCE", x"FD76", x"FD26", x"FCFD", x"FC43", x"FC0A", x"FC6A", x"FB4C", x"F8B9", x"F6A0", x"F546", x"F524", x"F7A4", x"FBDB", x"FF8D", x"02CB", x"05F0", x"0831", x"09EE", x"0BD7", x"0D15", x"0D2C", x"0CC5", x"0B8B", x"0980", x"0785", x"05B3", x"0393", x"01A6", x"FF9F", x"FCE0", x"F9E7", x"F74E", x"F45B", x"F176", x"EF5A", x"ED8F", x"EBF5", x"EB93", x"EBF4", x"EC56", x"ED73", x"EF5F", x"F10C", x"F313", x"F5BD", x"F7D3", x"F91C", x"FADB", x"FC92", x"FDC3", x"FF4C", x"006E", x"FF67", x"FD20", x"FB88", x"FAAE", x"FB78", x"FED0", x"0322", x"0696", x"09C9", x"0CE7", x"0F1C", x"10FD", x"12DD", x"13B7", x"1365", x"12D8", x"11BA", x"100A", x"0E99", x"0D4A", x"0BBB", x"0A5E", x"0927", x"0752", x"054B", x"0347", x"00AC", x"FDEA", x"FB9D", x"F982", x"F791", x"F692", x"F611", x"F5A6", x"F5FF", x"F6D3", x"F76B", x"F84E", x"F978", x"F9D3", x"F9CF", x"FA48", x"FAA4", x"FACC", x"FB92", x"FB7B", x"F935", x"F627", x"F3A3", x"F1C1", x"F1EE", x"F4D2", x"F859", x"FB65", x"FEB1", x"01D4", x"040B", x"0658", x"0896", x"0996", x"09AC", x"0987", x"085B", x"0691", x"0510", x"039C", x"021F", x"0176", x"011E", x"0068", x"FFBB", x"FEE6", x"FD41", x"FBAD", x"FAB7", x"FA0E", x"F9F6", x"FAFA", x"FC26", x"FD7D", x"FFAD", x"0226", x"0497", x"079B", x"0A76", x"0C06", x"0D0C", x"0DF2", x"0DE6", x"0DA9", x"0D9C", x"0BF5", x"0819", x"03E4", x"FFF5", x"FC90", x"FB71", x"FC72", x"FD7A", x"FE64", x"FFF1", x"0134", x"0200", x"0336", x"042B", x"0412", x"03B0", x"031A", x"01B4", x"0014", x"FEC1", x"FD52", x"FC08", x"FB70", x"FABF", x"F9C2", x"F8C8", x"F752", x"F520", x"F2F3", x"F0D3", x"EE87", x"EC9F", x"EB41", x"E9FC", x"E94C", x"E98A", x"E9FD", x"EAD5", x"EC70", x"EDC4", x"EE88", x"EF8E", x"F08D", x"F106", x"F203", x"F313", x"F26B", x"F087", x"EEE2", x"EDA0", x"ED9B", x"F04B", x"F482", x"F86E", x"FC5B", x"006D", x"0390", x"061C", x"08B4", x"0A3F", x"0A82", x"0A6E", x"09E1", x"086F", x"0706", x"05C4", x"042B", x"02B9", x"01EA", x"00F5", x"FFAB", x"FE57", x"FC4C", x"F95D", x"F680", x"F3D9", x"F128", x"EEF5", x"ED59", x"EC33", x"EC0A", x"ED3E", x"EF45", x"F21F", x"F578", x"F85D", x"FAA5", x"FCD5", x"FE8A", x"FFD4", x"016B", x"026D", x"017C", x"FF6B", x"FD43", x"FB38", x"FA8E", x"FC77", x"FF7C", x"0271", x"05CC", x"0903", x"0B05", x"0C6D", x"0D8A", x"0D76", x"0C91", x"0BC3", x"0A82", x"08AC", x"072C", x"05E7", x"0485", x"0402", x"041E", x"0414", x"03C2", x"030C", x"0111", x"FE20", x"FB49", x"F871", x"F5E6", x"F460", x"F35A", x"F2C5", x"F31A", x"F41C", x"F55D", x"F765", x"F9C8", x"FB5D", x"FCB3", x"FE3A", x"FF24", x"003E", x"0238", x"0344", x"0218", x"004E", x"FE6C", x"FC7D", x"FCA3", x"FF55", x"0249", x"04F6", x"0851", x"0B33", x"0CCB", x"0E51", x"0F35", x"0E64", x"0CF2", x"0BBA", x"09C4", x"07A4", x"061D", x"0493", x"0307", x"029B", x"02BB", x"02C3", x"02F4", x"02C2", x"0143", x"FF4A", x"FD7A", x"FB90", x"FA54", x"FA18", x"FA74", x"FB76", x"FD97", x"FFFC", x"0272", x"054B", x"0780", x"0861", x"08DB", x"08B6", x"079C", x"06DB", x"0691", x"04BC", x"0160", x"FDD0", x"F9EA", x"F687", x"F5A1", x"F69A", x"F7A8", x"F92C", x"FB45", x"FCC1", x"FDE7", x"FF64", x"0037", x"0029", x"0004", x"FF62", x"FE04", x"FCD6", x"FBE5", x"FAEC", x"FACA", x"FB8F", x"FC86", x"FDE6", x"FFA1", x"004A", x"FFC9", x"FEC5", x"FCEB", x"FA81", x"F8C0", x"F74D", x"F5C4", x"F4E2", x"F4A7", x"F441", x"F496", x"F5BC", x"F63D", x"F60F", x"F5F9", x"F511", x"F3E0", x"F420", x"F4F4", x"F46E", x"F33E", x"F1F6", x"F030", x"EFAB", x"F21B", x"F5E4", x"F9AC", x"FDFC", x"0215", x"04B2", x"06B2", x"0849", x"0870", x"07AF", x"06F9", x"059B", x"038F", x"0185", x"FF25", x"FC33", x"F9E3", x"F849", x"F6E9", x"F5FA", x"F54B", x"F3B5", x"F17A", x"EF5A", x"ED4F", x"EB8E", x"EAA8", x"EA67", x"EAB4", x"EBE8", x"EDD1", x"F003", x"F2D2", x"F5AF", x"F81E", x"FA70", x"FC87", x"FDCC", x"FF32", x"0169", x"030F", x"037C", x"0339", x"020C", x"0041", x"0008", x"01F3", x"04AB", x"07ED", x"0BC6", x"0EE0", x"10E8", x"129A", x"1387", x"1354", x"12E2", x"1244", x"10CE", x"0F44", x"0DBE", x"0BB1", x"09A7", x"0847", x"0706", x"0610", x"060C", x"05EA", x"04BF", x"0311", x"00D4", x"FDC8", x"FB25", x"F97C", x"F81F", x"F777", x"F7D5", x"F84D", x"F8F1", x"FA6E", x"FBCD", x"FC75", x"FD4E", x"FDF6", x"FDDA", x"FE65", x"FFBE", x"FFAF", x"FDD6", x"FB6C", x"F820", x"F4DF", x"F425", x"F5BF", x"F7DE", x"FAB4", x"FE7B", x"01AC", x"0412", x"0649", x"0775", x"0754", x"06EF", x"0658", x"0511", x"038D", x"0215", x"0057", x"FF47", x"FF29", x"FFA3", x"00AF", x"022B", x"02FA", x"02B6", x"01DA", x"005E", x"FEA4", x"FDB8", x"FDAF", x"FE47", x"0005", x"0292", x"053F", x"0852", x"0B8B", x"0DDB", x"0F60", x"106F", x"1051", x"0F82", x"0F8A", x"0FAB", x"0EA6", x"0CC1", x"0A03", x"0611", x"02AC", x"0190", x"01F2", x"033C", x"0596", x"0810", x"09BE", x"0B20", x"0C2D", x"0C87", x"0CBA", x"0CCB", x"0C19", x"0AC5", x"0931", x"06E4", x"0477", x"02CE", x"016E", x"005B", x"0080", x"0119", x"00C1", x"FF97", x"FD92", x"FA31", x"F672", x"F3AA", x"F150", x"EF71", x"EECD", x"EEEA", x"EF78", x"F119", x"F377", x"F557", x"F70D", x"F890", x"F903", x"F947", x"FA68", x"FB5B", x"FB22", x"FA7B", x"F942", x"F787", x"F755", x"F999", x"FD1B", x"0119", x"05DE", x"0A2D", x"0D50", x"0FC1", x"1155", x"11A6", x"114E", x"10DA", x"0FD4", x"0E53", x"0C80", x"0A2E", x"07AE", x"05AE", x"040B", x"02DD", x"023A", x"01A2", x"0037", x"FE1C", x"FB4B", x"F7D1", x"F457", x"F175", x"EF85", x"EEF2", x"EFF0", x"F1F5", x"F4C8", x"F80D", x"FB18", x"FDEE", x"00E9", x"0345", x"04C5", x"0674", x"085F", x"0953", x"095C", x"0891", x"0629", x"033B", x"020C", x"02BB", x"045B", x"06EB", x"09FC", x"0C0B", x"0D4D", x"0E44", x"0E68", x"0DD4", x"0D51", x"0CB8", x"0BA9", x"0A94", x"094A", x"0796", x"063C", x"0582", x"04FB", x"050B", x"05C6", x"05DA", x"04DA", x"030F", x"0019", x"FC55", x"F915", x"F6B1", x"F4CA", x"F408", x"F45D", x"F4EC", x"F618", x"F819", x"F9D4", x"FB3E", x"FCD7", x"FDCD", x"FE24", x"FF4C", x"0103", x"0176", x"00E0", x"FF8D", x"FCEA", x"FA6C", x"FA51", x"FC06", x"FE54", x"018F", x"055B", x"083C", x"0A4C", x"0BCE", x"0C34", x"0BA6", x"0B1B", x"0A87", x"0989", x"0829", x"066E", x"04C0", x"03D2", x"0394", x"0403", x"0549", x"06C0", x"0771", x"0770", x"065A", x"03D7", x"00E7", x"FED0", x"FD7E", x"FD52", x"FEB9", x"00D0", x"02F0", x"059A", x"083A", x"0A03", x"0B57", x"0C3B", x"0BCB", x"0AF7", x"0AFD", x"0AD9", x"09F0", x"088E", x"061F", x"025B", x"FF37", x"FDD1", x"FD52", x"FDCE", x"FF46", x"00B9", x"01C8", x"02F4", x"03F6", x"04AD", x"059C", x"065A", x"065D", x"0606", x"0540", x"03E0", x"02FD", x"02F8", x"02EC", x"037D", x"0571", x"0798", x"08F6", x"09B9", x"08F3", x"05ED", x"0257", x"FF4B", x"FC65", x"FA17", x"F931", x"F8F0", x"F921", x"FA5D", x"FBE9", x"FCF5", x"FDF9", x"FEC2", x"FEE5", x"FF3B", x"001B", x"009C", x"0075", x"0002", x"FEA5", x"FCEC", x"FC82", x"FDBA", x"0009", x"0370", x"0741", x"0A54", x"0C63", x"0DAD", x"0DEB", x"0DA3", x"0D46", x"0C7E", x"0B25", x"0978", x"0737", x"0493", x"028B", x"0100", x"FF74", x"FEAA", x"FEA3", x"FE64", x"FDAF", x"FC98", x"FA6F", x"F73B", x"F460", x"F21E", x"F074", x"F01E", x"F128", x"F303", x"F5B4", x"F909", x"FC1C", x"FF23", x"0246", x"04BD", x"06A8", x"08D8", x"0AD2", x"0BEE", x"0CA8", x"0C68", x"0A5A", x"07F6", x"06D9", x"06CA", x"07C9", x"0A1B", x"0C91", x"0E17", x"0F4F", x"103E", x"1041", x"0FF9", x"0FC6", x"0F09", x"0DEF", x"0CBC", x"0AFD", x"08DF", x"074B", x"0619", x"054E", x"05A0", x"06AD", x"0749", x"076B", x"06C4", x"04A2", x"01B3", x"FEFF", x"FC85", x"FA86", x"F9CA", x"F9C6", x"FA0C", x"FB07", x"FC2D", x"FCE6", x"FDD3", x"FECF", x"FEF1", x"FED8", x"FF56", x"FF75", x"FED5", x"FE1A", x"FC4A", x"F920", x"F6B9", x"F64B", x"F728", x"F962", x"FD1E", x"00CB", x"03E4", x"06E7", x"095A", x"0A75", x"0AC5", x"0A7C", x"0963", x"07DA", x"0619", x"0403", x"024B", x"0176", x"0123", x"01B2", x"0327", x"04A3", x"05CA", x"06B7", x"0698", x"050A", x"0340", x"01B0", x"0063", x"0065", x"01E2", x"03C3", x"0603", x"08E3", x"0B36", x"0CD0", x"0E61", x"0EF8", x"0E2A", x"0D61", x"0D13", x"0C50", x"0B7A", x"0A8C", x"07FD", x"0456", x"01C4", x"0092", x"0079", x"01ED", x"0461", x"063B", x"07E3", x"09A4", x"0ACD", x"0B80", x"0C06", x"0BF1", x"0AF7", x"098A", x"073B", x"0473", x"022D", x"0073", x"FF03", x"FE89", x"FEED", x"FF24", x"FF64", x"FF78", x"FE18", x"FB35", x"F800", x"F46F", x"F0DA", x"EE72", x"ED32", x"EC89", x"ED04", x"EE7D", x"EFFA", x"F17E", x"F336", x"F40B", x"F42F", x"F4B1", x"F535", x"F58D", x"F644", x"F6BF", x"F60A", x"F531", x"F58D", x"F6E2", x"F9A9", x"FE06", x"029E", x"0661", x"098D", x"0BB7", x"0CA8", x"0D01", x"0CF4", x"0BFD", x"0A90", x"08C4", x"063E", x"03C4", x"0201", x"005A", x"FEE4", x"FE3E", x"FDF3", x"FD74", x"FD3A", x"FCB8", x"FAD6", x"F82D", x"F596", x"F2FC", x"F0F7", x"F077", x"F10B", x"F262", x"F4E4", x"F7CB", x"FA76", x"FD15", x"FF85", x"0108", x"0244", x"038F", x"0458", x"049C", x"04C1", x"03BC", x"0140", x"FEC3", x"FD0C", x"FC39", x"FD19", x"FF96", x"0248", x"04A9", x"06DA", x"084E", x"08E9", x"093B", x"094F", x"08DB", x"0857", x"0793", x"0653", x"053D", x"0465", x"0380", x"02D7", x"02C2", x"0297", x"0255", x"0234", x"0160", x"FF75", x"FD29", x"FAC1", x"F84D", x"F6AD", x"F653", x"F6A8", x"F7DC", x"F9F6", x"FBEF", x"FDA7", x"FF72", x"00A7", x"00F2", x"013D", x"0190", x"014D", x"0118", x"00E5", x"FF3D", x"FC81", x"FA56", x"F927", x"F931", x"FB69", x"FF0C", x"0264", x"056B", x"084F", x"0A47", x"0B4B", x"0C00", x"0C04", x"0B35", x"0A2A", x"08DC", x"0733", x"05C1", x"04C4", x"03FE", x"03CD", x"041B", x"0457", x"046D", x"0454", x"0375", x"01C0", x"FFDA", x"FDE1", x"FC03", x"FB43", x"FB8E", x"FCA5", x"FEAA", x"0122", x"0311", x"0499", x"05D5", x"05F2", x"056B", x"04FD", x"0485", x"03C1", x"0370", x"02A2", x"FFF8", x"FC5E", x"F911", x"F650", x"F4DD", x"F57D", x"F700", x"F826", x"F98A", x"FB0F", x"FC26", x"FD17", x"FE28", x"FEC7", x"FEE8", x"FEEA", x"FE7C", x"FDAE", x"FD0F", x"FCA1", x"FC8F", x"FD10", x"FDD1", x"FE5E", x"FEE0", x"FEFD", x"FE0D", x"FC61", x"FA07", x"F6DF", x"F3B6", x"F176", x"EFFF", x"EF7A", x"F02F", x"F13D", x"F221", x"F347", x"F478", x"F4C0", x"F4ED", x"F55C", x"F592", x"F5E1", x"F703", x"F78B", x"F696", x"F587", x"F51E", x"F54C", x"F6FA", x"FA4B", x"FD6E", x"FF9D", x"0197", x"02E7", x"02FE", x"0285", x"01A3", x"000C", x"FE3F", x"FCC5", x"FB3D", x"F992", x"F82B", x"F6EF", x"F5FC", x"F596", x"F55D", x"F51A", x"F4C2", x"F415", x"F2A4", x"F0D9", x"EEB5", x"EC4E", x"EA68", x"E9A3", x"E9E0", x"EB5E", x"EE15", x"F130", x"F450", x"F7C8", x"FAED", x"FD66", x"FFDB", x"026B", x"0475", x"0684", x"085B", x"088E", x"06E6", x"04C0", x"02C4", x"0141", x"0169", x"02EB", x"0441", x"0552", x"0670", x"070B", x"06EF", x"06CF", x"069E", x"0631", x"05F5", x"05DE", x"0569", x"04DB", x"044D", x"03D5", x"03C3", x"0416", x"045D", x"049E", x"04CD", x"043A", x"02D1", x"00FA", x"FE90", x"FBC8", x"F9B2", x"F858", x"F76E", x"F76A", x"F839", x"F8E9", x"F9A2", x"FA96", x"FAB9", x"FA19", x"F9BE", x"F994", x"F94A", x"F9AC", x"FA0B", x"F8B2", x"F647", x"F445", x"F2D8", x"F2B8", x"F4E7", x"F82C", x"FACD", x"FD2B", x"FF4B", x"0037", x"0059", x"0053", x"FFA7", x"FE66", x"FD6B", x"FC9D", x"FBAC", x"FB31", x"FB50", x"FBB6", x"FCBE", x"FE49", x"FFC4", x"0121", x"0244", x"0286", x"01F3", x"00E1", x"FF46", x"FD84", x"FC7C", x"FC1B", x"FC7A", x"FDD1", x"FFAA", x"012F", x"02B4", x"03EC", x"0433", x"0432", x"0470", x"0470", x"047E", x"0518", x"050F", x"0368", x"015A", x"FF8D", x"FE30", x"FE77", x"00DA", x"037B", x"0597", x"07A7", x"0906", x"0974", x"09AB", x"09C8", x"090B", x"0804", x"06F4", x"0571", x"03AA", x"0226", x"00B1", x"FF6B", x"FEDF", x"FE97", x"FE69", x"FE8D", x"FE6C", x"FD7C", x"FC01", x"F9FB", x"F718", x"F463", x"F252", x"F0AD", x"EFDC", x"F027", x"F0A1", x"F118", x"F232", x"F31A", x"F33B", x"F377", x"F3E2", x"F3D5", x"F484", x"F62C", x"F71E", x"F6EA", x"F6DB", x"F6E3", x"F758", x"F9C1", x"FDC3", x"0154", x"0444", x"06EF", x"084F", x"0863", x"0814", x"071D", x"053E", x"0384", x"022A", x"00B3", x"FF4D", x"FE35", x"FD16", x"FC47", x"FBFF", x"FBE1", x"FBB4", x"FB89", x"FAD3", x"F9A5", x"F843", x"F684", x"F486", x"F307", x"F22C", x"F1ED", x"F309", x"F51A", x"F75D", x"F9F8", x"FCEE", x"FF29", x"00A8", x"0236", x"0334", x"03B8", x"04DA", x"0600", x"0569", x"0391", x"014B", x"FEAD", x"FCF9", x"FDB9", x"FFC5", x"01A8", x"038E", x"051E", x"0589", x"057B", x"058F", x"0538", x"0497", x"0459", x"0402", x"0360", x"02BB", x"0206", x"011C", x"0087", x"0031", x"FFD3", x"FFBB", x"FFB9", x"FF4B", x"FEA0", x"FDB8", x"FC2F", x"FA7B", x"F956", x"F885", x"F849", x"F92B", x"FA68", x"FB5C", x"FC9C", x"FDB9", x"FDAC", x"FD2F", x"FCA8", x"FB8A", x"FA79", x"FAB3", x"FAC1", x"F993", x"F806", x"F68B", x"F503", x"F54E", x"F813", x"FB93", x"FEC4", x"0217", x"04A8", x"05ED", x"06E8", x"07AE", x"076A", x"06D5", x"0671", x"05CA", x"04E8", x"0450", x"038E", x"029C", x"0200", x"01AD", x"0165", x"017F", x"01A7", x"0167", x"00CD", x"FFE6", x"FE65", x"FD03", x"FC1B", x"FBA8", x"FC11", x"FD6E", x"FED3", x"0025", x"01B7", x"02EB", x"036C", x"0403", x"0469", x"0405", x"03F1", x"047E", x"040F", x"0261", x"004C", x"FD91", x"FAE0", x"FA28", x"FB86", x"FD36", x"FF32", x"0161", x"02B9", x"0363", x"046D", x"054E", x"05B8", x"0647", x"06DD", x"06CD", x"0679", x"0606", x"051D", x"0434", x"03A5", x"031B", x"02AA", x"0268", x"01E9", x"00F1", x"FFDD", x"FE54", x"FC41", x"FA69", x"F8AB", x"F724", x"F692", x"F6D8", x"F745", x"F849", x"FA0B", x"FB59", x"FC3C", x"FD3B", x"FD8F", x"FD3E", x"FDD8", x"FF15", x"FF44", x"FEC8", x"FE05", x"FC7A", x"FB6B", x"FCAF", x"FF49", x"01B9", x"0438", x"063B", x"06AE", x"0668", x"0619", x"050F", x"0385", x"0264", x"0160", x"0032", x"FF77", x"FEFE", x"FE64", x"FE1A", x"FE2F", x"FE0F", x"FDEC", x"FDBE", x"FD10", x"FBF8", x"FAD3", x"F93B", x"F773", x"F5F4", x"F4BE", x"F420", x"F4D2", x"F68F", x"F8C8", x"FBEF", x"FF77", x"0272", x"053A", x"07F7", x"09E3", x"0B70", x"0DB3", x"0F64", x"0F70", x"0E4A", x"0C0B", x"08AB", x"0612", x"0593", x"05F5", x"068F", x"07AB", x"0860", x"0843", x"0846", x"0894", x"088D", x"088A", x"08FB", x"0919", x"0905", x"08F9", x"08BA", x"0832", x"07F0", x"07BE", x"078A", x"077E", x"0782", x"0709", x"0660", x"0552", x"03BE", x"01EF", x"0047", x"FE8C", x"FD60", x"FD10", x"FCF3", x"FD28", x"FDF5", x"FEA1", x"FEAE", x"FED4", x"FEA5", x"FD84", x"FCDD", x"FD2F", x"FD2F", x"FC81", x"FBC5", x"FA3D", x"F852", x"F83C", x"FA40", x"FCB8", x"FFA6", x"02B6", x"0499", x"0549", x"061A", x"067C", x"0610", x"05E3", x"0602", x"05C5", x"05A9", x"0612", x"0623", x"062D", x"06D3", x"07B9", x"089C", x"09D0", x"0AC8", x"0AD4", x"0A52", x"097A", x"0812", x"0684", x"0520", x"03CF", x"030B", x"0325", x"03BD", x"04D9", x"0660", x"07A0", x"087C", x"096C", x"09D3", x"09A1", x"09EB", x"0A91", x"0A6A", x"099B", x"0867", x"0645", x"043C", x"043B", x"05B9", x"077E", x"0997", x"0B64", x"0BCF", x"0B91", x"0B95", x"0B2D", x"0A5F", x"09E8", x"094C", x"0819", x"06E1", x"0599", x"03DE", x"0256", x"0170", x"00BA", x"0057", x"0042", x"FFE3", x"FF17", x"FE44", x"FD4C", x"FC15", x"FADE", x"F965", x"F7B4", x"F67E", x"F5AF", x"F524", x"F55F", x"F612", x"F688", x"F73F", x"F846", x"F8C3", x"F91A", x"FAB3", x"FC8D", x"FDD6", x"FF08", x"FFB6", x"FF31", x"FF4A", x"017C", x"044F", x"06FA", x"09C0", x"0B66", x"0B42", x"0AE0", x"0A84", x"0939", x"07A7", x"0693", x"054A", x"03FB", x"037F", x"0319", x"022D", x"019F", x"0156", x"00CE", x"0079", x"0059", x"FF83", x"FE2E", x"FD09", x"FBDF", x"FAB4", x"F9FD", x"F953", x"F8C1", x"F8CF", x"F981", x"FA8D", x"FC46", x"FE19", x"FF8A", x"00FD", x"0254", x"02EA", x"0398", x"0507", x"0614", x"0634", x"05CB", x"042D", x"017C", x"FFED", x"005A", x"0165", x"02FB", x"04F3", x"0610", x"063E", x"06E1", x"0789", x"07A1", x"07CC", x"0833", x"07F3", x"0796", x"0773", x"06D6", x"05F1", x"0588", x"0541", x"04FF", x"052D", x"0565", x"0521", x"04E3", x"04D0", x"0499", x"047B", x"047C", x"0424", x"03D9", x"03E1", x"03D4", x"03E9", x"046D", x"047E", x"042C", x"03FE", x"034D", x"01D7", x"013E", x"01B4", x"01DE", x"020F", x"0220", x"00F9", x"FF4D", x"FFB2", x"01B8", x"040F", x"0728", x"0A29", x"0B9C", x"0C55", x"0D98", x"0E39", x"0E20", x"0E63", x"0E76", x"0DB3", x"0D2E", x"0CB4", x"0B5B", x"09CF", x"08D9", x"07C8", x"06CB", x"0687", x"05FB", x"04CA", x"03BC", x"02D9", x"01D6", x"0132", x"00E5", x"005F", x"0016", x"005B", x"00D0", x"01B0", x"02EB", x"03B8", x"0425", x"0485", x"042B", x"0352", x"034B", x"0392", x"032E", x"0278", x"012D", x"FE69", x"FBF4", x"FB91", x"FC73", x"FDDD", x"0028", x"0212", x"02AD", x"0355", x"0467", x"04F2", x"0557", x"0631", x"0665", x"05F2", x"0594", x"04B7", x"031B", x"01C9", x"00E1", x"FFE3", x"FF71", x"FF78", x"FEF6", x"FE2D", x"FDA8", x"FCF9", x"FC56", x"FC31", x"FBD1", x"FB03", x"FA59", x"F9BD", x"F90E", x"F931", x"F9C5", x"FA10", x"FA85", x"FAFE", x"FA65", x"F9B3", x"FA2C", x"FAA4", x"FACD", x"FB2F", x"FAB9", x"F8FA", x"F836", x"F990", x"FB75", x"FDDE", x"00C3", x"0247", x"0241", x"026D", x"027B", x"0192", x"00CC", x"004D", x"FF31", x"FE2B", x"FDF6", x"FD6F", x"FC8F", x"FC3B", x"FBE0", x"FB37", x"FB13", x"FAF3", x"FA01", x"F8CC", x"F7CD", x"F6A4", x"F5E0", x"F5E5", x"F5EC", x"F61E", x"F6EE", x"F817", x"F9A9", x"FC24", x"FEBC", x"0117", x"039C", x"05A7", x"0683", x"077C", x"08CF", x"0965", x"096B", x"0914", x"06F1", x"0390", x"0175", x"00B3", x"0082", x"0175", x"02E6", x"032F", x"0315", x"03D6", x"047C", x"04D9", x"05D8", x"069F", x"0698", x"06B7", x"06FA", x"0679", x"05F9", x"05DF", x"0564", x"04DC", x"04C4", x"044C", x"031A", x"021D", x"0110", x"FFE1", x"FF3C", x"FEE2", x"FE1E", x"FD66", x"FCD3", x"FC0A", x"FB92", x"FBC6", x"FBAD", x"FB82", x"FB7D", x"FAAB", x"F911", x"F85C", x"F867", x"F84C", x"F8BF", x"F914", x"F7BF", x"F629", x"F639", x"F75E", x"F900", x"FBCA", x"FE39", x"FF11", x"FFA2", x"0089", x"00AD", x"00A2", x"0132", x"016C", x"015B", x"01DC", x"025E", x"0235", x"0248", x"02A2", x"02AD", x"02EC", x"0376", x"0334", x"0255", x"016D", x"003F", x"FF0C", x"FE71", x"FDFE", x"FD64", x"FD3D", x"FD5F", x"FDA3", x"FEB9", x"0039", x"0185", x"0304", x"0476", x"04DB", x"04DE", x"058D", x"060F", x"0642", x"06AA", x"0628", x"03EC", x"021E", x"01C2", x"020D", x"0333", x"054D", x"066E", x"0658", x"0682", x"06C4", x"0671", x"067B", x"06B5", x"0625", x"054A", x"04B8", x"037C", x"01E8", x"00C3", x"FF90", x"FE41", x"FDA4", x"FD47", x"FC63", x"FBA1", x"FAED", x"F9DF", x"F910", x"F8DD", x"F869", x"F7C1", x"F746", x"F66A", x"F565", x"F518", x"F4FD", x"F4E8", x"F559", x"F5D3", x"F570", x"F583", x"F689", x"F7AC", x"F91A", x"FAF7", x"FB9E", x"FAF7", x"FB18", x"FC37", x"FD8C", x"FF9D", x"01DE", x"028A", x"022E", x"01FF", x"0179", x"0082", x"0014", x"FFD0", x"FF1B", x"FEC7", x"FECB", x"FE62", x"FDF5", x"FDE4", x"FD9E", x"FD51", x"FD5E", x"FCFC", x"FC0E", x"FB0D", x"F9F4", x"F8E0", x"F861", x"F862", x"F84C", x"F862", x"F88F", x"F869", x"F89D", x"F946", x"F9F0", x"FAF5", x"FC80", x"FD8D", x"FDE7", x"FEBD", x"FF89", x"0005", x"00D0", x"0141", x"FFD8", x"FD92", x"FC28", x"FB48", x"FB31", x"FC87", x"FDEA", x"FE19", x"FE29", x"FE8B", x"FE8A", x"FEBA", x"FF98", x"001A", x"0021", x"0072", x"0076", x"FFF6", x"FFB4", x"FFB4", x"FF72", x"FF7E", x"FFCF", x"FFA3", x"FF24", x"FEC3", x"FE24", x"FD87", x"FD71", x"FD6E", x"FD06", x"FC8C", x"FBB6", x"FA68", x"F951", x"F897", x"F7BD", x"F741", x"F6FA", x"F610", x"F502", x"F4D0", x"F512", x"F5BD", x"F722", x"F821", x"F7AD", x"F713", x"F762", x"F833", x"F9C8", x"FC5F", x"FE67", x"FF5A", x"0029", x"00F1", x"0104", x"0126", x"0184", x"0179", x"014C", x"015C", x"0119", x"006E", x"FFE8", x"FF78", x"FEEC", x"FEC2", x"FE90", x"FDF2", x"FD1C", x"FC54", x"FB62", x"FAE2", x"FAFB", x"FB45", x"FBA3", x"FC36", x"FC7D", x"FC8E", x"FCED", x"FD3C", x"FD70", x"FDFC", x"FE5C", x"FDF1", x"FD82", x"FD75", x"FD3F", x"FD44", x"FDA8", x"FD04", x"FB24", x"F9A3", x"F902", x"F8F9", x"FA6F", x"FCC4", x"FE5F", x"FF2C", x"0004", x"0055", x"001C", x"003F", x"0062", x"FFED", x"FF8F", x"FF3D", x"FE57", x"FD4D", x"FCAB", x"FBF0", x"FB6F", x"FBA4", x"FBEC", x"FBD3", x"FBC6", x"FB88", x"FAD1", x"FA8D", x"FADE", x"FB26", x"FB64", x"FBA6", x"FB37", x"FA79", x"FA15", x"F9D4", x"F9AA", x"F9F5", x"F9FC", x"F94C", x"F8E5", x"F8EF", x"F923", x"F9FA", x"FB2D", x"FB3D", x"FA6B", x"FA07", x"F9F4", x"FA61", x"FBF8", x"FDE2", x"FEBF", x"FF2A", x"FF8F", x"FF39", x"FE9A", x"FE7E", x"FE2E", x"FDAE", x"FDA5", x"FDB8", x"FD3E", x"FCEE", x"FCC1", x"FC59", x"FC30", x"FC74", x"FC59", x"FBC8", x"FB38", x"FA42", x"F943", x"F901", x"F96A", x"F9FC", x"FAFE", x"FC00", x"FC93", x"FD28", x"FDF1", x"FE87", x"FF68", x"009F", x"0146", x"019B", x"022B", x"0292", x"02CB", x"0385", x"03C2", x"0270", x"00AD", x"FF52", x"FE19", x"FDDA", x"FF22", x"0039", x"008D", x"0115", x"0199", x"017B", x"01BC", x"025C", x"0250", x"0215", x"024A", x"022B", x"0192", x"015D", x"0100", x"002F", x"FFB7", x"FF75", x"FEAE", x"FDDF", x"FD29", x"FC1A", x"FB2E", x"FAF2", x"FAEE", x"FAE8", x"FB20", x"FB08", x"FA77", x"FA17", x"F9BA", x"F92E", x"F8FD", x"F8BF", x"F7D6", x"F6FF", x"F6BE", x"F6B3", x"F759", x"F8E7", x"F9D1", x"F973", x"F916", x"F8E3", x"F8D7", x"FA06", x"FC3A", x"FDC6", x"FEB0", x"FFD8", x"0084", x"00BD", x"0188", x"0261", x"02C5", x"035D", x"044A", x"04A9", x"04C3", x"0501", x"04D2", x"0469", x"045F", x"0424", x"0365", x"029A", x"0181", x"000A", x"FF08", x"FEB6", x"FEAB", x"FF3D", x"0028", x"00BA", x"011E", x"01C0", x"0218", x"0285", x"036B", x"0406", x"03E7", x"03F2", x"0419", x"0409", x"04BF", x"05DE", x"05E0", x"04DC", x"03FD", x"0309", x"0277", x"0384", x"0529", x"060F", x"069D", x"0706", x"067D", x"0594", x"051F", x"0458", x"0346", x"028F", x"01E6", x"00AA", x"FF88", x"FE8A", x"FD57", x"FC81", x"FC53", x"FC23", x"FBE0", x"FBBF", x"FB1C", x"FA39", x"F9B3", x"F98B", x"F983", x"FA0D", x"FA98", x"FA98", x"FA85", x"FA5B", x"F9E3", x"F9A4", x"F9DD", x"F9AE", x"F949", x"F95F", x"F98A", x"FA0C", x"FB9E", x"FD55", x"FDF4", x"FE0B", x"FE0E", x"FDBD", x"FE0D", x"FFA8", x"0134", x"01FB", x"02C3", x"0315", x"02BD", x"0293", x"02CD", x"02A5", x"0280", x"02D0", x"02D7", x"0296", x"0286", x"024F", x"01B5", x"016E", x"013A", x"0089", x"FFC5", x"FECB", x"FD58", x"FBF8", x"FB46", x"FAE4", x"FAF6", x"FB94", x"FC20", x"FC59", x"FCC2", x"FD06", x"FD19", x"FD8D", x"FE26", x"FE46", x"FE7B", x"FEE0", x"FF23", x"FF9F", x"00CB", x"0146", x"00A4", x"FFB3", x"FEA5", x"FD9A", x"FDE9", x"FF66", x"00A5", x"018F", x"0274", x"02CF", x"02AA", x"0303", x"0367", x"0356", x"0374", x"03C3", x"03A9", x"037C", x"038C", x"035F", x"0336", x"0381", x"03E9", x"0416", x"0457", x"044C", x"03D5", x"037A", x"0363", x"0366", x"03B0", x"0424", x"0433", x"0406", x"03BB", x"030A", x"0253", x"01FE", x"0179", x"00C9", x"006E", x"003C", x"0035", x"0137", x"02E3", x"03D6", x"0405", x"03D7", x"02E6", x"0221", x"02AD", x"03F9", x"04EB", x"05F2", x"06E5", x"070B", x"071D", x"0793", x"07C3", x"07AB", x"0802", x"0864", x"085A", x"0865", x"0843", x"079B", x"06D2", x"0659", x"05A9", x"04E3", x"0418", x"02F3", x"0187", x"0080", x"FFF7", x"FFFC", x"00D0", x"01F3", x"02FC", x"03DF", x"0466", x"045E", x"044F", x"0450", x"03F7", x"038E", x"034F", x"02D3", x"027A", x"02F3", x"0389", x"0349", x"02C2", x"01DD", x"009F", x"0018", x"0104", x"0232", x"030B", x"03D7", x"0403", x"036B", x"02EB", x"02CE", x"0266", x"0213", x"021C", x"01F2", x"0187", x"0140", x"00EF", x"0080", x"0078", x"00C3", x"00FA", x"0128", x"0118", x"00A2", x"0003", x"FFA2", x"FF60", x"FF89", x"0006", x"007A", x"00DF", x"0130", x"00F8", x"0051", x"FFB0", x"FED6", x"FD9D", x"FCB0", x"FC08", x"FB49", x"FB70", x"FCA0", x"FDB4", x"FE28", x"FE58", x"FDC3", x"FCBC", x"FCB5", x"FDC9", x"FEC1", x"FF9F", x"0079", x"0090", x"003D", x"0069", x"00B3", x"00BC", x"00F9", x"017A", x"0196", x"01AB", x"01DB", x"01AF", x"0165", x"014D", x"0128", x"00C0", x"0037", x"FF59", x"FE26", x"FD45", x"FCDD", x"FD03", x"FDE1", x"FF31", x"006B", x"01A4", x"02A9", x"030A", x"0346", x"03A2", x"03D2", x"03F0", x"045C", x"0497", x"046A", x"04D8", x"059E", x"05C7", x"0582", x"04FC", x"03BB", x"028B", x"029C", x"035F", x"0404", x"04C4", x"054F", x"0519", x"04C2", x"04CB", x"04A3", x"0465", x"048B", x"04C8", x"04E8", x"052F", x"055E", x"052A", x"04FD", x"04D1", x"0495", x"044A", x"0404", x"0342", x"0255", x"016C", x"0077", x"FFCF", x"FFC6", x"FFEA", x"0032", x"00A5", x"00BD", x"002E", x"FFA3", x"FF13", x"FE31", x"FDA2", x"FD72", x"FD16", x"FD05", x"FE16", x"FF6E", x"005C", x"011C", x"0126", x"003B", x"FFA6", x"002E", x"011B", x"021C", x"0365", x"0424", x"043A", x"0467", x"04BF", x"04B9", x"04C5", x"04FC", x"04F0", x"04C0", x"04C3", x"049C", x"047A", x"048E", x"04A9", x"0478", x"0435", x"0395", x"0297", x"01B0", x"00F7", x"0085", x"0099", x"013C", x"01F2", x"02E5", x"03D4", x"0445", x"0442", x"044B", x"0403", x"039B", x"0399", x"03AE", x"0383", x"03E3", x"04FB", x"05DD", x"067A", x"06D2", x"0639", x"050D", x"04AC", x"053F", x"060D", x"071B", x"0803", x"07F1", x"0747", x"06CE", x"0669", x"05FF", x"0604", x"05F6", x"057C", x"04B6", x"03D5", x"02B5", x"01DE", x"0181", x"015B", x"0143", x"0124", x"009E", x"FFCA", x"FEFA", x"FE3A", x"FDAE", x"FDA2", x"FDDB", x"FE42", x"FEEF", x"FF94", x"FFCA", x"FFCE", x"FFAD", x"FF22", x"FE9D", x"FE70", x"FE2D", x"FDDF", x"FE61", x"FF56", x"0035", x"0109", x"018B", x"00F3", x"FFF3", x"FF9E", x"FFAA", x"FFF3", x"009C", x"0148", x"014D", x"0147", x"0185", x"01A7", x"01C2", x"0238", x"028A", x"02A5", x"0299", x"025A", x"01B8", x"0118", x"009B", x"001F", x"FFA0", x"FF0E", x"FE2D", x"FD30", x"FC63", x"FBD1", x"FBC9", x"FC52", x"FD17", x"FE08", x"FF0B", x"FF9F", x"FF96", x"FF66", x"FEF6", x"FE5B", x"FE34", x"FE7A", x"FE7B", x"FE91", x"FF36", x"FFE0", x"005E", x"010F", x"0150", x"00C3", x"0060", x"00CD", x"0160", x"0221", x"031B", x"0383", x"0342", x"031A", x"032F", x"0329", x"0370", x"0411", x"0484", x"04D1", x"0520", x"0515", x"04AF", x"0452", x"03E7", x"0358", x"02DD", x"0246", x"016B", x"0091", x"FFCD", x"FF27", x"FEE3", x"FF0B", x"FF43", x"FFAB", x"0021", x"002C", x"FFDC", x"FF8D", x"FEE4", x"FE1E", x"FDBC", x"FD7D", x"FD0C", x"FD1E", x"FDE6", x"FEBB", x"FF82", x"0037", x"FFDD", x"FEA3", x"FDBB", x"FD7A", x"FD99", x"FE49", x"FF3E", x"FF9A", x"FF8D", x"FFB6", x"FFE0", x"0012", x"00AA", x"0149", x"01A8", x"01E5", x"01F7", x"01C9", x"01A9", x"01BC", x"01AC", x"0180", x"011B", x"0039", x"FF25", x"FE3C", x"FD82", x"FD32", x"FD96", x"FE4E", x"FF43", x"0084", x"01AF", x"0235", x"026A", x"0251", x"018F", x"00D5", x"007C", x"FFE6", x"FF30", x"FF0E", x"FF3D", x"FF6A", x"FFEF", x"0069", x"FFEA", x"FF16", x"FECC", x"FED8", x"FF2F", x"FFFA", x"0088", x"0034", x"FFAF", x"FF41", x"FEC5", x"FE90", x"FED0", x"FF0C", x"FF34", x"FF6C", x"FF79", x"FF68", x"FF94", x"FFE0", x"0033", x"0081", x"00A6", x"0048", x"FFB3", x"FEF4", x"FE05", x"FD3C", x"FCCF", x"FC8D", x"FCB1", x"FD46", x"FDC4", x"FDF4", x"FDF9", x"FD75", x"FC7B", x"FBB3", x"FB33", x"FA95", x"FA3E", x"FA7B", x"FABE", x"FB0B", x"FB92", x"FB94", x"FAA9", x"F9AD", x"F90D", x"F8A7", x"F8D5", x"F98F", x"FA21", x"FA70", x"FAFF", x"FBB1", x"FC7C", x"FD8C", x"FED0", x"FFD5", x"00B1", x"0153", x"018A", x"0184", x"0183", x"0165", x"013C", x"0112", x"0090", x"FFCC", x"FF03", x"FE39", x"FD9F", x"FD78", x"FDB1", x"FE05", x"FEA1", x"FF53", x"FFA3", x"FFC5", x"FFD1", x"FF8B", x"FF34", x"FF4A", x"FF65", x"FF3E", x"FF58", x"FFB8", x"FFF9", x"0077", x"012D", x"012F", x"009D", x"002D", x"0008", x"0010", x"00AC", x"0160", x"016E", x"00FD", x"0086", x"FFE6", x"FF76", x"FF7C", x"FFC5", x"FFE9", x"001D", x"0017", x"FFBD", x"FF58", x"FF0E", x"FEBD", x"FE73", x"FE3C", x"FDA7", x"FCEF", x"FC25", x"FB53", x"FA9E", x"FA53", x"FA3F", x"FA4F", x"FAA7", x"FAF7", x"FAF3", x"FAD8", x"FA9B", x"FA00", x"F993", x"F98C", x"F97F", x"F987", x"FA10", x"FADB", x"FBAD", x"FCE7", x"FDF7", x"FE18", x"FDAE", x"FD52", x"FD04", x"FD19", x"FDE8", x"FEB9", x"FF12", x"FF50", x"FF7C", x"FF84", x"FFC1", x"0055", x"00B8", x"00FE", x"0136", x"0139", x"010B", x"0104", x"00F8", x"00AE", x"004F", x"FFB3", x"FECC", x"FDDD", x"FD33", x"FCAA", x"FC8E", x"FCE0", x"FD5F", x"FE04", x"FEEC", x"FFA1", x"0027", x"007F", x"005C", x"FFB0", x"FF1B", x"FE9B", x"FE1C", x"FDEE", x"FE51", x"FEC2", x"FF73", x"008A", x"014A", x"014B", x"0115", x"00CA", x"0071", x"0074", x"00D6", x"00DA", x"006A", x"FFDE", x"FF36", x"FE82", x"FE3D", x"FE2C", x"FE12", x"FDF1", x"FDCA", x"FD59", x"FCF4", x"FCB4", x"FC91", x"FC81", x"FC90", x"FC62", x"FBF1", x"FB57", x"FAAB", x"F9F6", x"F9A3", x"F985", x"F9A0", x"FA0B", x"FAAB", x"FB34", x"FBB6", x"FC0C", x"FBBD", x"FB1A", x"FA84", x"F9E3", x"F93B", x"F922", x"F95E", x"F9C9", x"FAA2", x"FBE4", x"FC8E", x"FC85", x"FC49", x"FBE8", x"FB8D", x"FBE9", x"FCA8", x"FD19", x"FD3E", x"FD6D", x"FD7C", x"FD8C", x"FE07", x"FE9D", x"FEF5", x"FF3A", x"FF40", x"FEDB", x"FE2B", x"FD75", x"FCB0", x"FBF0", x"FB55", x"FAA1", x"F9B7", x"F8C3", x"F7DF", x"F73B", x"F720", x"F772", x"F80B", x"F8D1", x"F974", x"F9EA", x"FA3B", x"FA6F", x"FA57", x"FA42", x"FA41", x"FA13", x"F9C3", x"F9BA", x"F9CE", x"FA13", x"FAED", x"FC0A", x"FCA8", x"FCD2", x"FCE8", x"FCCA", x"FCD0", x"FD5B", x"FDF1", x"FDFF", x"FDD1", x"FDA5", x"FD68", x"FD7D", x"FE25", x"FEF4", x"FFB6", x"0071", x"00F5", x"010A", x"010F", x"00FD", x"00CE", x"00A7", x"006C", x"0003", x"FF70", x"FEF5", x"FE5E", x"FE05", x"FDEA", x"FDED", x"FE16", x"FE7F", x"FEEA", x"FF27", x"FF69", x"FF6B", x"FF02", x"FEB7", x"FE8A", x"FE31", x"FDEF", x"FE1E", x"FE5B", x"FED0", x"FFDB", x"00C7", x"00E5", x"00A5", x"0045", x"FFAE", x"FF85", x"0016", x"008B", x"0097", x"00AB", x"00A2", x"0075", x"00A7", x"0126", x"015B", x"015B", x"015B", x"0101", x"008E", x"0065", x"0040", x"0009", x"FFE9", x"FFAE", x"FF39", x"FED6", x"FEA1", x"FE79", x"FE9C", x"FF07", x"FF7C", x"000E", x"00BE", x"0146", x"019C", x"01E4", x"01A6", x"0114", x"0070", x"FFBC", x"FEC2", x"FE11", x"FDAE", x"FD60", x"FD97", x"FE60", x"FED3", x"FEC1", x"FE63", x"FDB1", x"FCD2", x"FC8F", x"FCBC", x"FCB4", x"FC77", x"FC33", x"FBAA", x"FB4F", x"FB94", x"FC38", x"FCFA", x"FDF4", x"FEB8", x"FF21", x"FF65", x"FFAC", x"FFCE", x"0002", x"004A", x"004C", x"0007", x"FFAA", x"FF00", x"FE3D", x"FDBE", x"FD6A", x"FD3E", x"FD70", x"FDC3", x"FDEE", x"FE19", x"FE17", x"FD92", x"FCD3", x"FC2A", x"FB37", x"FA3B", x"F99C", x"F934", x"F8F0", x"F97C", x"FA68", x"FAF7", x"FB0D", x"FAE6", x"FA4E", x"F9AC", x"F9DF", x"FA56", x"FAAD", x"FB05", x"FB64", x"FB99", x"FC1E", x"FD2A", x"FE4B", x"FF3E", x"001D", x"0084", x"007C", x"0051", x"0023", x"FFE0", x"FFBF", x"FFB7", x"FF7F", x"FF39", x"FEF7", x"FEAA", x"FE82", x"FEAA", x"FEF5", x"FF57", x"FFDF", x"004A", x"008D", x"00D2", x"00F8", x"00D6", x"00BA", x"0095", x"001E", x"FF96", x"FF4C", x"FF0C", x"FF1D", x"FFFD", x"00F8", x"018F", x"01C9", x"01B6", x"0133", x"00F7", x"0169", x"01CE", x"01E4", x"01C9", x"0167", x"00C1", x"0094", x"00DB", x"0143", x"01B0", x"023E", x"025F", x"0262", x"0256", x"023F", x"01F7", x"01D6", x"0181", x"00F6", x"0060", x"FFC5", x"FF06", x"FE79", x"FE30", x"FDE9", x"FDD9", x"FE17", x"FE47", x"FE7E", x"FEE8", x"FF25", x"FF2F", x"FF59", x"FF6C", x"FF13", x"FEC9", x"FEB5", x"FE94", x"FF05", x"0032", x"0156", x"01F6", x"0259", x"022D", x"0190", x"0164", x"01C3", x"01F6", x"0211", x"0225", x"01DB", x"0179", x"0199", x"01F1", x"0233", x"0293", x"02CC", x"029A", x"024F", x"0215", x"01BD", x"017F", x"017C", x"0152", x"0119", x"00F9", x"00C8", x"009E", x"00B9", x"00F1", x"0125", x"01A4", x"0241", x"02C1", x"034E", x"03CD", x"03C0", x"0377", x"033A", x"029E", x"01E3", x"016E", x"0127", x"0107", x"01CD", x"032A", x"043F", x"0500", x"0561", x"0505", x"048A", x"04A9", x"051B", x"055A", x"0599", x"0598", x"051D", x"04D9", x"0508", x"0559", x"05B8", x"0639", x"0660", x"0619", x"05D0", x"0552", x"04BE", x"0450", x"0402", x"0384", x"0303", x"0277", x"01BA", x"010F", x"00B7", x"006F", x"0065", x"00A5", x"00E6", x"0115", x"0161", x"0192", x"0178", x"0176", x"0174", x"0115", x"00A0", x"0044", x"FFCA", x"FF84", x"FFFB", x"00B0", x"011E", x"0151", x"0128", x"0072", x"FFEA", x"0002", x"0047", x"0092", x"00EB", x"011A", x"011A", x"016E", x"021F", x"02EC", x"03BC", x"0473", x"049F", x"0451", x"03BE", x"02F4", x"0223", x"018B", x"0107", x"006A", x"FFE2", x"FF4A", x"FEB0", x"FE5C", x"FE4B", x"FE50", x"FE90", x"FEF2", x"FF39", x"FF73", x"FFBF", x"FFDA", x"FFD7", x"FFFB", x"000D", x"FFC9", x"FF82", x"FF4E", x"FF21", x"FF7F", x"00D9", x"025D", x"03AC", x"04A8", x"0500", x"04AA", x"048B", x"04D8", x"052B", x"0561", x"05A4", x"0583", x"0529", x"0535", x"0583", x"05E3", x"0678", x"0710", x"0746", x"0745", x"0728", x"06C8", x"0652", x"0600", x"0589", x"04F8", x"0471", x"03DC", x"032C", x"02B6", x"026C", x"0234", x"023B", x"028E", x"02BD", x"02F5", x"0340", x"034D", x"0341", x"035A", x"033A", x"02CD", x"0263", x"0207", x"01A6", x"01E0", x"02A9", x"0354", x"03B0", x"03BA", x"0330", x"0244", x"01E1", x"01E1", x"01EB", x"0220", x"0257", x"0238", x"021E", x"0275", x"02E4", x"036D", x"041E", x"0497", x"04A2", x"0482", x"043B", x"03BD", x"0373", x"0359", x"0340", x"0336", x"0351", x"0341", x"0327", x"033A", x"033C", x"0340", x"038F", x"03F4", x"044E", x"04DC", x"0557", x"057E", x"0583", x"0578", x"04DC", x"0415", x"0357", x"028D", x"01FA", x"0244", x"0300", x"03A2", x"0420", x"042C", x"0365", x"0276", x"01FA", x"019B", x"013C", x"010E", x"0091", x"FFCC", x"FF58", x"FF6E", x"FFC4", x"0084", x"0193", x"024C", x"02C1", x"0310", x"0313", x"02E6", x"02E2", x"02FA", x"02E9", x"02E1", x"02A6", x"021E", x"017B", x"0106", x"00A7", x"0092", x"00D3", x"0113", x"0140", x"016F", x"015A", x"010F", x"00D3", x"0084", x"FFE8", x"FF3D", x"FE84", x"FD99", x"FCFB", x"FD17", x"FD7B", x"FDE1", x"FE46", x"FE3D", x"FDBB", x"FD6A", x"FDA7", x"FE0E", x"FEB8", x"FF80", x"001D", x"0087", x"0143", x"0233", x"0335", x"0454", x"056D", x"0622", x"0677", x"068A", x"063C", x"05B6", x"054C", x"04DE", x"0464", x"03FD", x"0386", x"0301", x"02AC", x"0287", x"0288", x"02AF", x"02E3", x"02F3", x"0302", x"0317", x"0314", x"0310", x"0336", x"032A", x"02DB", x"0283", x"0201", x"0177", x"016C", x"021D", x"02F7", x"03C0", x"045B", x"0437", x"038F", x"031A", x"02F0", x"02D1", x"02D7", x"02D4", x"027B", x"01F5", x"01C2", x"01AD", x"01B9", x"0212", x"025E", x"0265", x"0242", x"01FB", x"016F", x"00FF", x"00B1", x"0052", x"FFE7", x"FF89", x"FEFB", x"FE5A", x"FDF9", x"FDB2", x"FD88", x"FDAD", x"FE01", x"FE40", x"FE97", x"FEFF", x"FF18", x"FF41", x"FF7D", x"FF7D", x"FF40", x"FF0B", x"FEB4", x"FE65", x"FEE0", x"FFFC", x"012C", x"023D", x"02F4", x"02C6", x"022D", x"01E1", x"01D7", x"01D5", x"0228", x"0268", x"024C", x"0236", x"025A", x"027B", x"02B4", x"032F", x"037E", x"0395", x"0388", x"0343", x"02B1", x"0241", x"01FA", x"01AF", x"0190", x"017A", x"012D", x"00D8", x"009C", x"0070", x"006E", x"00BE", x"0118", x"016F", x"01D5", x"020A", x"0206", x"01FC", x"01D8", x"0166", x"00DE", x"005D", x"FFAD", x"FF4E", x"FFA5", x"0063", x"0139", x"022D", x"0297", x"024D", x"01DB", x"0196", x"015B", x"0159", x"0186", x"0179", x"0131", x"0121", x"0136", x"0188", x"0240", x"0326", x"03BD", x"0422", x"042A", x"03CB", x"0345", x"02E5", x"0272", x"0207", x"01A6", x"0115", x"005C", x"FFB6", x"FF2D", x"FEA4", x"FE72", x"FE69", x"FE50", x"FE52", x"FE60", x"FE2D", x"FDED", x"FDEA", x"FDCC", x"FD8C", x"FD5A", x"FCF6", x"FC32", x"FBC5", x"FBFB", x"FC62", x"FCFC", x"FD9F", x"FDAF", x"FD32", x"FCE2", x"FCEE", x"FD1C", x"FD9C", x"FE54", x"FEAF", x"FEF3", x"FF5F", x"FFDC", x"005A", x"0100", x"0181", x"01A4", x"0169", x"00F1", x"001D", x"FF3B", x"FE7D", x"FDC3", x"FD0B", x"FC56", x"FB8B", x"FAB1", x"FA1B", x"F9C4", x"F9C5", x"FA14", x"FA70", x"FAC1", x"FB1A", x"FB5D", x"FB95", x"FBE5", x"FC4C", x"FC7B", x"FC8E", x"FC8D", x"FC41", x"FBF8", x"FC2E", x"FCF5", x"FDF5", x"FF2B", x"001F", x"0056", x"0006", x"FFBB", x"FF7E", x"FF76", x"FFC1", x"0010", x"0011", x"FFF3", x"FFC2", x"FF9E", x"FFBA", x"0031", x"00A6", x"0112", x"0143", x"0117", x"00B7", x"006F", x"0013", x"FFB6", x"FF5E", x"FEED", x"FE45", x"FDBB", x"FD5C", x"FD13", x"FD11", x"FD72", x"FDD0", x"FE3A", x"FEC6", x"FF1C", x"FF2A", x"FF64", x"FF92", x"FF91", x"FF95", x"FF9B", x"FF17", x"FEA0", x"FE9B", x"FEF5", x"FF7C", x"0048", x"00BD", x"0053", x"FFA5", x"FF17", x"FE8F", x"FE59", x"FE8D", x"FEB4", x"FEA1", x"FEA9", x"FEBD", x"FECB", x"FF0D", x"FF86", x"FFD1", x"000B", x"0025", x"FFF9", x"FFA8", x"FF7F", x"FF69", x"FF7C", x"FFC2", x"0012", x"0034", x"0052", x"005D", x"005E", x"007F", x"00B1", x"00D7", x"00FB", x"0124", x"011B", x"010A", x"00F6", x"00A5", x"0016", x"FF85", x"FEB9", x"FDC2", x"FD25", x"FD05", x"FD3A", x"FDC7", x"FE7A", x"FE97", x"FE1C", x"FD76", x"FCC3", x"FC26", x"FBF2", x"FBE0", x"FBA3", x"FB4D", x"FB1D", x"FAFF", x"FB50", x"FC1E", x"FD15", x"FE09", x"FED5", x"FF3D", x"FF45", x"FF48", x"FF3B", x"FF17", x"FEEA", x"FEA2", x"FDE9", x"FD29", x"FC7A", x"FBDD", x"FB7B", x"FB82", x"FB89", x"FB87", x"FBAA", x"FBA4", x"FB54", x"FB17", x"FAF4", x"FA9C", x"FA60", x"FA42", x"F9BB", x"F8DD", x"F854", x"F812", x"F80D", x"F888", x"F922", x"F91B", x"F8B8", x"F879", x"F84C", x"F86A", x"F913", x"F9DD", x"FA61", x"FAE1", x"FB71", x"FBED", x"FC9E", x"FD88", x"FE6B", x"FF28", x"FFBC", x"FFFF", x"FFE4", x"FFB5", x"FF71", x"FF18", x"FECC", x"FE7E", x"FE02", x"FD9F", x"FD40", x"FD01", x"FCF1", x"FD10", x"FD24", x"FD3D", x"FD60", x"FD67", x"FD56", x"FD78", x"FD95", x"FD92", x"FDB8", x"FDC6", x"FD74", x"FD15", x"FD0C", x"FD2D", x"FDAB", x"FE7E", x"FF26", x"FF27", x"FEDD", x"FE75", x"FDFC", x"FDC4", x"FDEC", x"FE0A", x"FE13", x"FE16", x"FDF9", x"FDEC", x"FE07", x"FE5F", x"FEA5", x"FEFA", x"FF13", x"FEDC", x"FEA3", x"FE63", x"FE1C", x"FDD1", x"FD8B", x"FCFF", x"FC55", x"FBD6", x"FB66", x"FB22", x"FB4A", x"FBA0", x"FBEB", x"FC68", x"FCE8", x"FD2C", x"FD64", x"FDC3", x"FDEE", x"FDFE", x"FE48", x"FE4B", x"FDEB", x"FD9F", x"FD9C", x"FDAD", x"FE30", x"FEF4", x"FF48", x"FEED", x"FE68", x"FDCA", x"FD31", x"FD31", x"FD78", x"FDB1", x"FDBD", x"FDCA", x"FDA1", x"FD8F", x"FDC2", x"FE1C", x"FE6C", x"FEC0", x"FED7", x"FEA4", x"FE6F", x"FE33", x"FDFA", x"FDD9", x"FDBF", x"FD87", x"FD31", x"FCFA", x"FCB2", x"FC8E", x"FCA9", x"FCC5", x"FCE3", x"FD0B", x"FD28", x"FD13", x"FD28", x"FD4F", x"FD5C", x"FD77", x"FDA6", x"FD83", x"FD32", x"FD10", x"FD27", x"FD70", x"FE42", x"FF25", x"FF9D", x"FFA5", x"FF7D", x"FF30", x"FEFF", x"FF3A", x"FF8F", x"FFC1", x"FFE6", x"FFEA", x"FFED", x"0021", x"00A0", x"014D", x"0206", x"02A3", x"02DF", x"02C4", x"0277", x"01FE", x"017F", x"0114", x"0079", x"FFBF", x"FEEF", x"FE2D", x"FD6A", x"FD08", x"FCE4", x"FCC9", x"FCD2", x"FCED", x"FCD3", x"FCAC", x"FC9D", x"FC81", x"FC57", x"FC6F", x"FC95", x"FC70", x"FC44", x"FC28", x"FC02", x"FC08", x"FC76", x"FCD3", x"FCB7", x"FC76", x"FC00", x"FB82", x"FB4B", x"FB9D", x"FC04", x"FC6E", x"FCD8", x"FD28", x"FD47", x"FD90", x"FDE0", x"FE3F", x"FE93", x"FEE5", x"FEF1", x"FECA", x"FE7F", x"FE0A", x"FD86", x"FCF8", x"FC56", x"FB99", x"FAEB", x"FA54", x"F9F1", x"F9E4", x"FA13", x"FA54", x"FAB6", x"FB14", x"FB52", x"FB9E", x"FBFF", x"FC64", x"FCCE", x"FD6B", x"FDE8", x"FE2E", x"FE75", x"FED7", x"FF4D", x"0003", x"00FB", x"01AD", x"01DD", x"01C4", x"0180", x"012A", x"0117", x"0158", x"018C", x"01A0", x"01A4", x"0192", x"0162", x"0154", x"017B", x"01B7", x"01FE", x"0240", x"0253", x"022A", x"01DF", x"0195", x"0153", x"00FE", x"009B", x"000A", x"FF65", x"FEC9", x"FE87", x"FE9C", x"FEE0", x"FF49", x"FFB4", x"FFF2", x"000F", x"003B", x"006F", x"0088", x"00C4", x"010D", x"010D", x"00E2", x"00A7", x"0076", x"0050", x"0091", x"0102", x"0116", x"00C5", x"0036", x"FF69", x"FEBD", x"FE75", x"FE9A", x"FEBE", x"FEF0", x"FF1F", x"FF2C", x"FF21", x"FF3E", x"FF77", x"FFCA", x"003A", x"00AE", x"00F9", x"0130", x"0151", x"0184", x"01CD", x"0216", x"025A", x"0285", x"029A", x"02A6", x"02BE", x"02EC", x"0313", x"032F", x"0347", x"0337", x"0304", x"02DB", x"02A2", x"0262", x"0233", x"0210", x"01C4", x"0158", x"0107", x"00D7", x"00C3", x"0110", x"0162", x"015E", x"00FE", x"0082", x"FFE6", x"FF58", x"FF29", x"FF18", x"FEFE", x"FEE2", x"FEE9", x"FEED", x"FEF8", x"FF47", x"FFC9", x"006A", x"0126", x"01E0", x"0251", x"0279", x"0285", x"027E", x"0263", x"0238", x"01F2", x"0187", x"0113", x"00C7", x"00B2", x"00C6", x"00EC", x"0117", x"0119", x"00ED", x"00BA", x"007A", x"003E", x"000F", x"FFFB", x"FFDC", x"FF94", x"FF46", x"FEEF", x"FE99", x"FE79", x"FE9B", x"FEB8", x"FEA1", x"FE71", x"FE24", x"FDE7", x"FE00", x"FE93", x"FF4F", x"0023", x"00F4", x"01AA", x"022A", x"02B1", x"0340", x"03E1", x"0487", x"0530", x"05AD", x"05D5", x"05C4", x"058D", x"053B", x"04E8", x"0483", x"040E", x"0377", x"02F3", x"0284", x"0258", x"024C", x"0266", x"0282", x"0285", x"0279", x"026D", x"0272", x"0290", x"02C2", x"0308", x"0328", x"0323", x"0307", x"02EF", x"02E6", x"031C", x"0385", x"03C7", x"03BF", x"0384", x"031D", x"02B0", x"0282", x"02A0", x"02C3", x"02DA", x"02F4", x"02EC", x"02B4", x"0287", x"027E", x"0285", x"029C", x"02E6", x"0305", x"02E5", x"02A3", x"0270", x"0220", x"01DE", x"0194", x"0126", x"0086", x"0015", x"FFF3", x"0016", x"007C", x"0111", x"0184", x"01D2", x"0217", x"025B", x"029C", x"02E0", x"0341", x"0387", x"03AF", x"03BA", x"03BF", x"03A8", x"03B0", x"03E7", x"0423", x"0432", x"03FD", x"0399", x"0317", x"02AC", x"0296", x"02C9", x"0305", x"0344", x"037A", x"037F", x"0350", x"0331", x"0323", x"0338", x"036D", x"03CB", x"0403", x"03F5", x"03D6", x"03AC", x"0376", x"0347", x"031E", x"02C8", x"0263", x"0211", x"01F2", x"01E4", x"01FF", x"0217", x"0210", x"01F3", x"01D8", x"01CD", x"01D4", x"01FA", x"022B", x"0250", x"025D", x"024E", x"0242", x"0243", x"026D", x"02C2", x"0328", x"0360", x"035E", x"0346", x"0316", x"02F5", x"0314", x"0371", x"03CF", x"043F", x"04C2", x"0516", x"0547", x"058D", x"05F3", x"0665", x"06FC", x"079A", x"07D8", x"07B8", x"076E", x"0702", x"0675", x"05EF", x"055A", x"0483", x"03A5", x"02DF", x"0251", x"01E2", x"01C6", x"01A1", x"0173", x"0139", x"0107", x"00D7", x"00D0", x"00F0", x"0120", x"014E", x"0178", x"0185", x"0188", x"0190", x"01A7", x"01C4", x"01D3", x"01AE", x"0155", x"00D7", x"0058", x"0006", x"0007", x"004E", x"00AE", x"011E", x"0185", x"01AC", x"01B4", x"01C2", x"01DE", x"020E", x"0275", x"02DC", x"02E9", x"02BF", x"0262", x"01CD", x"012A", x"008F", x"FFE1", x"FF09", x"FE55", x"FDCB", x"FD6F", x"FD5D", x"FD78", x"FD92", x"FDA0", x"FDC5", x"FDFA", x"FE54", x"FEE5", x"FF91", x"002C", x"00B8", x"012F", x"017D", x"01D7", x"023B", x"02A9", x"031D", x"0372", x"0397", x"0379", x"0340", x"02F2", x"02BD", x"02BB", x"02BD", x"02C2", x"02C5", x"02B3", x"026E", x"022E", x"0200", x"01D5", x"01CE", x"0207", x"022D", x"022C", x"0224", x"0217", x"01F5", x"01DC", x"01D5", x"0195", x"0138", x"00FF", x"00F5", x"010E", x"016B", x"01CF", x"020F", x"0229", x"0246", x"0253", x"0276", x"02AE", x"02FE", x"0332", x"0362", x"0373", x"036B", x"0360", x"035A", x"035F", x"035C", x"0331", x"02CF", x"0245", x"019F", x"0110", x"00B7", x"00A8", x"00AD", x"00CC", x"00FC", x"0103", x"00DC", x"00C2", x"00A6", x"00B0", x"0104", x"01AB", x"0247", x"02C2", x"0340", x"0397", x"03DC", x"042D", x"0476", x"047B", x"045A", x"0441", x"041B", x"03FD", x"03FA", x"03E9", x"03A8", x"035E", x"0309", x"02A3", x"0248", x"0207", x"01B9", x"0171", x"011E", x"00C9", x"006A", x"0024", x"FFFC", x"FFE6", x"FFEC", x"FFE1", x"FFB5", x"FF6B", x"FF0D", x"FEAD", x"FE75", x"FE6E", x"FE70", x"FE94", x"FEC8", x"FEDD", x"FEDA", x"FEE2", x"FF01", x"FF2C", x"FFAC", x"0042", x"00AD", x"00E9", x"010A", x"00FA", x"00CF", x"00AC", x"006B", x"FFF8", x"FF79", x"FF13", x"FEAE", x"FE78", x"FE63", x"FE54", x"FE34", x"FE1A", x"FDF2", x"FDCF", x"FDC1", x"FDCB", x"FDCF", x"FDCE", x"FDCC", x"FDA5", x"FD8A", x"FD77", x"FD78", x"FD7C", x"FD8A", x"FD70", x"FD37", x"FCF0", x"FCAA", x"FC9A", x"FCD6", x"FD4A", x"FDD4", x"FE82", x"FF14", x"FF79", x"FFBA", x"FFF6", x"0015", x"004C", x"00B2", x"0115", x"013E", x"0155", x"0142", x"0109", x"00CB", x"009F", x"0047", x"FFCE", x"FF6A", x"FF07", x"FEB6", x"FEA7", x"FEAA", x"FEAF", x"FEC2", x"FEE3", x"FF0B", x"FF4E", x"FFAF", x"000D", x"0051", x"0074", x"007F", x"0059", x"003D", x"002B", x"0029", x"0032", x"0045", x"002D", x"0004", x"FFB3", x"FF66", x"FF38", x"FF35", x"FF44", x"FF68", x"FF9A", x"FFB2", x"FFAD", x"FFA3", x"FF87", x"FF5A", x"FF56", x"FF84", x"FFA1", x"FFAF", x"FFB0", x"FF8A", x"FF4A", x"FF18", x"FEE8", x"FE9C", x"FE51", x"FE22", x"FE00", x"FE08", x"FE46", x"FE90", x"FEE3", x"FF2B", x"FF7E", x"FFB2", x"FFF1", x"002B", x"0056", x"006D", x"0084", x"0079", x"006B", x"004A", x"002A", x"0006", x"FFE4", x"FFA7", x"FF53", x"FEE1", x"FE58", x"FDE2", x"FDAA", x"FD9D", x"FDAF", x"FDF1", x"FE3E", x"FE76", x"FEA1", x"FEC5", x"FECE", x"FEDE", x"FF29", x"FF98", x"FFF2", x"003E", x"005E", x"0046", x"000F", x"FFDB", x"FF9A", x"FF37", x"FECB", x"FE58", x"FDD7", x"FD65", x"FD0F", x"FCBD", x"FC7F", x"FC53", x"FC3E", x"FC33", x"FC44", x"FC68", x"FC93", x"FCCB", x"FD05", x"FD40", x"FD6F", x"FDA1", x"FDE1", x"FE39", x"FE94", x"FEDE", x"FF0C", x"FEFD", x"FED8", x"FEC6", x"FEE1", x"FF19", x"FF6E", x"FFF0", x"0066", x"00CC", x"012E", x"0176", x"01A6", x"01E5", x"0250", x"02B9", x"02F7", x"0316", x"02EB", x"0289", x"0210", x"0192", x"00F6", x"003A", x"FF84", x"FEC4", x"FE1E", x"FDA3", x"FD52", x"FD13", x"FCF2", x"FCD6", x"FCD2", x"FCCD", x"FCEA", x"FD09", x"FD26", x"FD45", x"FD61", x"FD73", x"FD70", x"FD78", x"FD7F", x"FD91", x"FD97", x"FD79", x"FD37", x"FCAA", x"FC2B", x"FBC8", x"FBA6", x"FBA9", x"FBDE", x"FC3C", x"FC88", x"FCD0", x"FD11", x"FD32", x"FD39", x"FD61", x"FDA5", x"FDE9", x"FE14", x"FE28", x"FE04", x"FDBB", x"FD5E", x"FCFD", x"FC6C", x"FBE2", x"FB46", x"FABA", x"FA3D", x"F9E6", x"F9B4", x"F9A1", x"F9C5", x"FA0C", x"FA80", x"FB11", x"FBBF", x"FC68", x"FD07", x"FD8C", x"FDF2", x"FE49", x"FE81", x"FEB9", x"FF04", x"FF48", x"FF74", x"FF8B", x"FF68", x"FF11", x"FEB1", x"FE80", x"FE48", x"FE22", x"FE19", x"FE1E", x"FE0F", x"FE04", x"FDFA", x"FDB3", x"FD70", x"FD4F", x"FD5D", x"FD71", x"FD98", x"FDBC", x"FDB7", x"FDAB", x"FDA9", x"FD9A", x"FD7C", x"FD58", x"FD31", x"FD00", x"FCE2", x"FCD7", x"FCDC", x"FCE9", x"FD05", x"FD27", x"FD4D", x"FD7E", x"FDB6", x"FDE8", x"FE11", x"FE36", x"FE51", x"FE57", x"FE4B", x"FE3C", x"FE31", x"FE1B", x"FE01", x"FDD7", x"FD70", x"FCEF", x"FC84", x"FC37", x"FC07", x"FC02", x"FC1A", x"FC2E", x"FC33", x"FC4D", x"FC53", x"FC53", x"FC70", x"FCC2", x"FD36", x"FDBE", x"FE51", x"FECA", x"FF2A", x"FF86", x"FFE2", x"002F", x"0066", x"0078", x"0058", x"001F", x"FFD1", x"FF87", x"FF46", x"FF0B", x"FED1", x"FE9C", x"FE64", x"FE39", x"FE0F", x"FDF5", x"FDD6", x"FDBC", x"FDA1", x"FD6C", x"FD3A", x"FD1D", x"FD21", x"FD2E", x"FD51", x"FD4E", x"FD1C", x"FCC5", x"FC92", x"FC73", x"FC65", x"FC85", x"FCB5", x"FCCC", x"FCE5", x"FCF8", x"FCF8", x"FCDE", x"FCF0", x"FD30", x"FD7A", x"FDCB", x"FE0D", x"FE1C", x"FDFA", x"FDE2", x"FDC2", x"FD91", x"FD4E", x"FD03", x"FCAE", x"FC5A", x"FC44", x"FC40", x"FC51", x"FC64", x"FC84", x"FC95", x"FCA2", x"FCBD", x"FCC5", x"FCC0", x"FCB6", x"FCC5", x"FCC2", x"FCB6", x"FCAF", x"FCBC", x"FCC1", x"FCE0", x"FCF3", x"FCE1", x"FC8D", x"FC4B", x"FC28", x"FC28", x"FC59", x"FCC8", x"FD3F", x"FDBA", x"FE30", x"FEAA", x"FEDF", x"FF03", x"FF32", x"FF5E", x"FF8F", x"FFBF", x"FFDA", x"FFCB", x"FFA0", x"FF7E", x"FF4F", x"FF10", x"FECD", x"FE78", x"FE17", x"FDC4", x"FD98", x"FD89", x"FD9E", x"FDD3", x"FE28", x"FE89", x"FEF5", x"FF64", x"FFB6", x"FFF0", x"000A", x"0010", x"FFFB", x"FFCC", x"FFAA", x"FFA2", x"FFA2", x"FFB0", x"FFAF", x"FF7F", x"FF1A", x"FEBE", x"FE84", x"FE4A", x"FE34", x"FE3D", x"FE4D", x"FE4B", x"FE5C", x"FE60", x"FE2D", x"FE0E", x"FE02", x"FE29", x"FE41", x"FE7A", x"FE9B", x"FE93", x"FE8E", x"FE95", x"FE95", x"FE79", x"FE52", x"FE18", x"FDC6", x"FD97", x"FD8E", x"FDAA", x"FDD7", x"FE2C", x"FE7F", x"FED8", x"FF20", x"FF6E", x"FF97", x"FFB3", x"FFD7", x"FFED", x"FFF0", x"FFD9", x"FFDB", x"FFCF", x"FFD6", x"FFF4", x"FFF6", x"FFB2", x"FF58", x"FEF8", x"FEBA", x"FE94", x"FEBF", x"FEEF", x"FF2A", x"FF5B", x"FFA0", x"FFC2", x"FFE4", x"0016", x"005D", x"009F", x"00E2", x"0117", x"0117", x"00FF", x"00E9", x"00D5", x"00C1", x"009A", x"0061", x"FFFC", x"FF81", x"FF11", x"FEB5", x"FE69", x"FE3A", x"FE24", x"FE18", x"FE18", x"FE36", x"FE58", x"FE84", x"FEBB", x"FF0B", x"FF48", x"FF85", x"FFB1", x"FFE2", x"000C", x"0049", x"0097", x"00BD", x"00C5", x"00BA", x"00BA", x"00D9", x"0118", x"0193", x"020C", x"028B", x"02F0", x"0358", x"038D", x"03BA", x"03F3", x"0441", x"0487", x"04BA", x"04D8", x"04A7", x"044C", x"03F1", x"0392", x"0306", x"0266", x"01BC", x"00EC", x"002C", x"FFAF", x"FF52", x"FF03", x"FEDC", x"FED8", x"FED4", x"FEE9", x"FF20", x"FF48", x"FF4E", x"FF7B", x"FFA4", x"FFCB", x"FFED", x"001F", x"0031", x"0044", x"006C", x"0084", x"006B", x"001B", x"FFCB", x"FF6D", x"FF37", x"FF37", x"FF66", x"FF9C", x"FFD2", x"000A", x"002E", x"0026", x"0013", x"001A", x"0025", x"004A", x"0084", x"00BA", x"00BD", x"00B8", x"00B8", x"009F", x"005E", x"000D", x"FF8A", x"FEE0", x"FE54", x"FDF9", x"FDC3", x"FDB9", x"FDF0", x"FE37", x"FE99", x"FF1F", x"FFB6", x"0032", x"00AD", x"0123", x"018A", x"01E5", x"0246", x"029E", x"02F1", x"0342", x"0398", x"03C2", x"03B9", x"037A", x"032A", x"02D7", x"029F", x"0288", x"0287", x"0283", x"0260", x"0243", x"01F8", x"0193", x"012C", x"00FD", x"00DB", x"00E0", x"0107", x"012A", x"0138", x"015F", x"01AA", x"01DE", x"020F", x"0224", x"0213", x"01D8", x"01B5", x"01B0", x"01AC", x"01BF", x"01F7", x"022B", x"0268", x"02BF", x"0305", x"0326", x"0339", x"0350", x"0351", x"0346", x"0349", x"033F", x"032A", x"0330", x"034D", x"0340", x"0301", x"029A", x"0227", x"01A8", x"016A", x"0169", x"0169", x"0179", x"019A", x"01BD", x"01E1", x"0208", x"0257", x"02B4", x"0326", x"03B3", x"0444", x"04BC", x"0518", x"0584", x"05D8", x"061B", x"0634", x"0622", x"05CF", x"0553", x"04E6", x"047A", x"0415", x"03C2", x"0385", x"0342", x"0314", x"02FF", x"02E2", x"02A9", x"0284", x"0261", x"0238", x"0227", x"021C", x"0207", x"01E2", x"01EF", x"01FA", x"01ED", x"01D8", x"01AC", x"0179", x"0152", x"0162", x"0188", x"01AF", x"01CF", x"01F2", x"01FD", x"01FD", x"01FE", x"0215", x"0242", x"0278", x"02AF", x"02D4", x"02C7", x"0295", x"026D", x"023E", x"01EC", x"0199", x"013A", x"00C1", x"0060", x"0033", x"001D", x"0003", x"000A", x"0016", x"0014", x"0031", x"0062", x"0078", x"0074", x"009B", x"00B7", x"00DD", x"011C", x"015A", x"0163", x"0176", x"0199", x"01A9", x"0190", x"0163", x"0115", x"00AA", x"006E", x"006D", x"008A", x"00CB", x"011E", x"0178", x"01BB", x"01EE", x"0208", x"0223", x"0236", x"025D", x"0284", x"02AE", x"02BB", x"02CA", x"02DA", x"02DF", x"02C2", x"029E", x"024E", x"01EA", x"0196", x"0171", x"0166", x"0185", x"01D0", x"0223", x"0277", x"02E4", x"033C", x"0365", x"0378", x"0383", x"0376", x"0374", x"0389", x"0394", x"0384", x"0390", x"03A0", x"039F", x"037D", x"0350", x"02F7", x"029D", x"0268", x"0263", x"0267", x"0275", x"028B", x"0289", x"0271", x"024C", x"0227", x"0212", x"020C", x"022F", x"0266", x"02A6", x"02E4", x"032B", x"0380", x"03B5", x"03DF", x"03E0", x"03B0", x"0359", x"030D", x"02C4", x"028B", x"0267", x"026B", x"027A", x"02A4", x"02FD", x"0347", x"0364", x"0385", x"0391", x"038A", x"0388", x"03A2", x"0386", x"0356", x"0342", x"032E", x"02F7", x"02AA", x"0248", x"01A9", x"0116", x"00C5", x"00A5", x"00A3", x"00C7", x"010C", x"0145", x"0190", x"01E1", x"0237", x"027A", x"02CB", x"0303", x"0337", x"0355", x"0361", x"0371", x"0377", x"036E", x"033B", x"02F4", x"0272", x"01CD", x"0133", x"0092", x"FFF4", x"FF71", x"FF1E", x"FED6", x"FECC", x"FEEF", x"FF1A", x"FF33", x"FF70", x"FFBB", x"0006", x"0078", x"00F0", x"0139", x"0174", x"01CB", x"021C", x"0252", x"0292", x"02B8", x"02B9", x"02D1", x"030D", x"0358", x"03A2", x"03F7", x"0437", x"0462", x"047F", x"0498", x"04AF", x"04D8", x"0501", x"0527", x"053D", x"0528", x"04F8", x"04C2", x"0479", x"0410", x"0396", x"0307", x"024D", x"019A", x"010C", x"0080", x"0011", x"FFCF", x"FFA6", x"FF8C", x"FFAA", x"FFDD", x"FFF3", x"000E", x"0032", x"0052", x"006F", x"00BA", x"00D9", x"00DD", x"00D7", x"00D8", x"00C2", x"00A7", x"0086", x"0037", x"FFC6", x"FF7D", x"FF3B", x"FF22", x"FF23", x"FF3C", x"FF38", x"FF2C", x"FF19", x"FEF2", x"FEEE", x"FEEF", x"FF0F", x"FF26", x"FF52", x"FF67", x"FF7B", x"FF8C", x"FF98", x"FF7B", x"FF5E", x"FF15", x"FEB7", x"FE5F", x"FE1F", x"FE00", x"FE0E", x"FE4F", x"FEAA", x"FF0F", x"FF87", x"FFEA", x"002C", x"0060", x"0095", x"00BC", x"00F9", x"014F", x"0186", x"01B7", x"01EB", x"0221", x"0243", x"0251", x"0242", x"01EC", x"0182", x"0120", x"00DC", x"00A4", x"008D", x"0075", x"004B", x"000D", x"FFD0", x"FF8A", x"FF53", x"FF2A", x"FF2F", x"FF36", x"FF5A", x"FF7A", x"FFA6", x"FFC3", x"FFE9", x"0001", x"000E", x"FFEE", x"FFBB", x"FF7A", x"FF41", x"FF0B", x"FF01", x"FF04", x"FF0B", x"FF35", x"FF6C", x"FF91", x"FFA1", x"FFA9", x"FFA2", x"FF8C", x"FF9B", x"FFBC", x"FFBE", x"FFCE", x"FFEF", x"0014", x"002B", x"003A", x"0020", x"FFB5", x"FF40", x"FEE7", x"FE98", x"FE76", x"FE84", x"FE9B", x"FEBA", x"FEE9", x"FF27", x"FF68", x"FFB9", x"0029", x"0091", x"010A", x"0173", x"01CE", x"0216", x"0250", x"0270", x"0273", x"025D", x"0216", x"01BA", x"015A", x"00EE", x"0077", x"0017", x"FFBC", x"FF70", x"FF46", x"FF42", x"FF29", x"FF0D", x"FEFD", x"FEE8", x"FECD", x"FECA", x"FEBC", x"FE8E", x"FE5F", x"FE5B", x"FE59", x"FE5C", x"FE66", x"FE51", x"FE0F", x"FDDE", x"FDBF", x"FDB1", x"FDBB", x"FDD3", x"FDE3", x"FDE2", x"FDDC", x"FDCF", x"FDC6", x"FDD1", x"FDE4", x"FE09", x"FE1B", x"FE11", x"FDF3", x"FDCF", x"FDA8", x"FD85", x"FD70", x"FD4E", x"FD17", x"FCF4", x"FCD5", x"FCBF", x"FCBD", x"FCDD", x"FCFA", x"FD22", x"FD67", x"FDA4", x"FDD2", x"FE06", x"FE48", x"FE77", x"FEB0", x"FEE0", x"FEEA", x"FECD", x"FEB0", x"FE87", x"FE58", x"FE39", x"FE02", x"FDBC", x"FD5B", x"FD13", x"FCDF", x"FCD9", x"FD0C", x"FD4E", x"FD98", x"FDCB", x"FDF1", x"FDF8", x"FE13", x"FE36", x"FE6E", x"FEA9", x"FEE3", x"FF06", x"FF23", x"FF3D", x"FF4F", x"FF5A", x"FF54", x"FF2E", x"FEEB", x"FE9B", x"FE4B", x"FE07", x"FDE6", x"FDE1", x"FDFF", x"FE16", x"FE46", x"FE55", x"FE5D", x"FE66", x"FE69", x"FE76", x"FE79", x"FE7A", x"FE60", x"FE33", x"FE19", x"FDFB", x"FDFA", x"FDFC", x"FDFA", x"FDD8", x"FDA4", x"FD72", x"FD47", x"FD2E", x"FD32", x"FD33", x"FD28", x"FD0F", x"FCEF", x"FCC4", x"FC9B", x"FC94", x"FC99", x"FCC9", x"FD0B", x"FD67", x"FDBE", x"FE13", x"FE59", x"FE8F", x"FE9E", x"FE8F", x"FE55", x"FE03", x"FDAC", x"FD55", x"FD27", x"FD0B", x"FD0B", x"FD1E", x"FD51", x"FD74", x"FDB2", x"FDE7", x"FE1E", x"FE42", x"FE6A", x"FE7C", x"FE77", x"FE67", x"FE6B", x"FE64", x"FE6A", x"FE66", x"FE41", x"FDD7", x"FD6D", x"FCF7", x"FC9A", x"FC68", x"FC69", x"FC7D", x"FC9D", x"FCD4", x"FD06", x"FD39", x"FD75", x"FDB8", x"FDFA", x"FE3D", x"FE7A", x"FE9F", x"FEB7", x"FEBF", x"FEB7", x"FE9F", x"FE76", x"FE27", x"FDC2", x"FD52", x"FCCD", x"FC48", x"FBE3", x"FB7E", x"FB44", x"FB27", x"FB3E", x"FB4B", x"FB81", x"FBBF", x"FC05", x"FC4E", x"FCAB", x"FCEC", x"FD1B", x"FD54", x"FDA2", x"FDFE", x"FE81", x"FF00", x"FF56", x"FF85", x"FFA4", x"FFAD", x"FFC2", x"FFE6", x"0010", x"0029", x"003D", x"0040", x"003F", x"0042", x"005E", x"0085", x"00B9", x"00DE", x"00DD", x"00BA", x"0082", x"002A", x"FFCC", x"FF70", x"FEFF", x"FE82", x"FE06", x"FD88", x"FD0C", x"FCA6", x"FC6C", x"FC3D", x"FC40", x"FC55", x"FC7C", x"FC98", x"FCC7", x"FCE9", x"FD0D", x"FD34", x"FD51", x"FD5D", x"FD51", x"FD55", x"FD44", x"FD53", x"FD66", x"FD75", x"FD63", x"FD4E", x"FD17", x"FCE6", x"FCAF", x"FC97", x"FC70", x"FC5B", x"FC3B", x"FC19", x"FBF7", x"FBEA", x"FBED", x"FC06", x"FC31", x"FC50", x"FC69", x"FC7B", x"FC97", x"FCA8", x"FCC6", x"FCDE", x"FCDF", x"FCD6", x"FCC7", x"FCB3", x"FC9D", x"FC9A", x"FCA1", x"FCAB", x"FCBF", x"FCD8", x"FCE4", x"FCFC", x"FD16", x"FD33", x"FD54", x"FD89", x"FDB8", x"FDE0", x"FE18", x"FE4A", x"FE8B", x"FED5", x"FF2F", x"FF6B", x"FF7E", x"FF7D", x"FF51", x"FF1C", x"FEF2", x"FECD", x"FEA4", x"FE6C", x"FE32", x"FDD9", x"FD7C", x"FD2D", x"FCE4", x"FCBB", x"FCAC", x"FCB5", x"FCD1", x"FCFB", x"FD37", x"FD66", x"FD93", x"FDB9", x"FDCB", x"FDD3", x"FDD5", x"FDD5", x"FDC5", x"FDCD", x"FDD5", x"FDE3", x"FDFE", x"FE22", x"FE3A", x"FE6C", x"FE94", x"FEC6", x"FEEB", x"FF1A", x"FF2B", x"FF36", x"FF43", x"FF56", x"FF79", x"FFB6", x"FFFA", x"0014", x"0015", x"FFED", x"FFB0", x"FF7E", x"FF73", x"FF84", x"FFAE", x"FFE5", x"0013", x"002B", x"0048", x"0060", x"0085", x"00C6", x"010B", x"0152", x"018A", x"01CF", x"01F4", x"0212", x"022A", x"0224", x"01FB", x"01D3", x"0189", x"0127", x"00A7", x"002D", x"FF99", x"FF24", x"FEDB", x"FEAF", x"FEA2", x"FEBE", x"FED2", x"FEDD", x"FEE4", x"FEE6", x"FEC8", x"FEAD", x"FE9E", x"FE7C", x"FE7E", x"FE98", x"FEB4", x"FEBA", x"FEC0", x"FEAE", x"FE8E", x"FE8E", x"FEA5", x"FEC3", x"FEEA", x"FF0E", x"FF05", x"FEF5", x"FEE8", x"FEDD", x"FED0", x"FEDA", x"FEC9", x"FE9C", x"FE6F", x"FE47", x"FE0C", x"FDDD", x"FDB8", x"FD80", x"FD56", x"FD43", x"FD38", x"FD31", x"FD35", x"FD43", x"FD4F", x"FD79", x"FDB3", x"FDFB", x"FE5E", x"FEC2", x"FF14", x"FF53", x"FF80", x"FF87", x"FF81", x"FF7B", x"FF62", x"FF40", x"FF2D", x"FF21", x"FF09", x"FF04", x"FEF8", x"FEDC", x"FEC3", x"FEC3", x"FEC1", x"FED7", x"FF00", x"FF20", x"FF2E", x"FF47", x"FF67", x"FF85", x"FFC3", x"FFFE", x"0027", x"003D", x"0065", x"007E", x"0099", x"00BF", x"00D4", x"00D2", x"00C3", x"00B2", x"0090", x"007A", x"006F", x"0067", x"0066", x"0073", x"007B", x"008C", x"00BB", x"00E3", x"0100", x"0120", x"0129", x"011B", x"0110", x"0102", x"00EA", x"00D7", x"00F3", x"0117", x"0148", x"0173", x"018B", x"0174", x"0162", x"014F", x"0142", x"0143", x"0143", x"0134", x"0108", x"00E9", x"00C2", x"00BC", x"00D3", x"0112", x"0144", x"0199", x"01E1", x"022C", x"025D", x"0284", x"0288", x"0267", x"023B", x"0200", x"01BB", x"0184", x"0150", x"012D", x"0119", x"0112", x"0120", x"0139", x"017E", x"01B7", x"01F6", x"0225", x"0231", x"022C", x"0218", x"020B", x"01F4", x"01FB", x"020D", x"021E", x"0215", x"01F1", x"0198", x"012F", x"00CD", x"0081", x"005E", x"0066", x"0094", x"00B6", x"00EF", x"012A", x"015E", x"01B2", x"0219", x"026F", x"02A9", x"02D9", x"02F5", x"02F3", x"02F1", x"02DF", x"029D", x"0240", x"01EA", x"0176", x"0100", x"0085", x"0000", x"FF72", x"FF03", x"FEBC", x"FEA6", x"FECB", x"FF20", x"FF85", x"FFE7", x"004D", x"0090", x"00DA", x"012A", x"018F", x"01FC", x"0286", x"030E", x"0385", x"03E8", x"042C", x"0441", x"0449", x"0450", x"0445", x"044F", x"045D", x"045F", x"0443", x"0433", x"0413", x"0404", x"0415", x"0444", x"0452", x"0446", x"0437", x"0407", x"03C6", x"039E", x"035E", x"031A", x"02CE", x"0295", x"0250", x"0203", x"01BC", x"0172", x"0131", x"0114", x"0108", x"0123", x"014D", x"0194", x"01CE", x"0216", x"022D", x"0237", x"0230", x"022D", x"021B", x"021F", x"0224", x"0223", x"0229", x"0232", x"0222", x"01F6", x"01C7", x"0185", x"0141", x"0124", x"011D", x"0103", x"00F0", x"00DB", x"00B9", x"00B0", x"00D1", x"0104", x"0126", x"0154", x"017A", x"0198", x"01C3", x"0205", x"0240", x"0275", x"02A5", x"02C9", x"02CE", x"02BD", x"0293", x"025D", x"0227", x"01F6", x"01CB", x"01B7", x"01AD", x"01BB", x"01DE", x"0202", x"0221", x"0234", x"0253", x"026B", x"0294", x"02D1", x"0314", x"035A", x"039F", x"03D2", x"03E0", x"03D2", x"03B4", x"0385", x"035A", x"033D", x"0317", x"02DB", x"029B", x"0247", x"01F0", x"01B0", x"0194", x"018B", x"0192", x"01B1", x"01DD", x"0209", x"0240", x"0276", x"0296", x"02A8", x"02B6", x"02C1", x"02B3", x"02AA", x"0289", x"0270", x"0245", x"022D", x"021F", x"0222", x"0243", x"0274", x"02B1", x"02D9", x"02EA", x"02E4", x"02CF", x"02C6", x"02D7", x"0309", x"034A", x"039D", x"03DA", x"0401", x"0403", x"03FB", x"03E0", x"03C7", x"03BE", x"03C8", x"03C9", x"03D2", x"03C9", x"03BA", x"03AC", x"03B6", x"03E5", x"0409", x"043A", x"046A", x"048E", x"04A0", x"04C1", x"04CF", x"04C2", x"04A5", x"0488", x"0451", x"03FD", x"0399", x"0319", x"0290", x"0215", x"01C5", x"0195", x"018B", x"01A8", x"01D1", x"01FC", x"021A", x"0223", x"0209", x"01E7", x"01C1", x"01B0", x"01AF", x"01C2", x"01E0", x"01F1", x"01F9", x"01ED", x"01E8", x"01D5", x"01D7", x"01DF", x"01F7", x"01FD", x"01FC", x"01E3", x"01BB", x"018C", x"0190", x"0197", x"019F", x"01A4", x"0193", x"0168", x"0131", x"0106", x"00DD", x"00AF", x"009C", x"00AC", x"00B3", x"00CC", x"00DE", x"00F1", x"0100", x"012F", x"0177", x"01C5", x"021A", x"026E", x"02B8", x"02E6", x"02FB", x"02F0", x"02C4", x"0285", x"0250", x"021D", x"0205", x"01F4", x"01EC", x"01D8", x"01BD", x"0198", x"0179", x"0153", x"013B", x"0131", x"0126", x"0117", x"0108", x"00FD", x"00E2", x"00F6", x"0126", x"016B", x"01A5", x"01E4", x"020B", x"021D", x"0231", x"024D", x"0255", x"024D", x"0257", x"0257", x"024A", x"023A", x"0220", x"01EE", x"01BD", x"019F", x"0190", x"017F", x"018C", x"0198", x"01B1", x"01BD", x"01C8", x"01B4", x"019B", x"0179", x"016F", x"0172", x"0199", x"01C0", x"01E6", x"01F9", x"01FA", x"01E7", x"01D6", x"01BD", x"01B2", x"01AC", x"0197", x"017B", x"0157", x"0124", x"00FE", x"00F0", x"010F", x"0136", x"015F", x"0194", x"01AA", x"01BC", x"01C7", x"01D5", x"01B7", x"0189", x"0163", x"011E", x"00DA", x"008A", x"0042", x"FFDF", x"FFA0", x"FF79", x"FF6D", x"FF6F", x"FF95", x"FFC9", x"0006", x"0050", x"008F", x"00B5", x"00C7", x"00D5", x"00DE", x"00FD", x"0124", x"014A", x"0155", x"0139", x"00FC", x"0099", x"003B", x"FFE0", x"FFA7", x"FF8B", x"FF76", x"FF6D", x"FF5C", x"FF4E", x"FF47", x"FF74", x"FFB9", x"000D", x"005D", x"00A7", x"00C7", x"00CE", x"00E1", x"00D4", x"00B5", x"008F", x"0069", x"0026", x"FFD2", x"FF7F", x"FF03", x"FE80", x"FE16", x"FDD0", x"FDA5", x"FDAD", x"FDE2", x"FE26", x"FE90", x"FEFA", x"FF67", x"FFB8", x"0008", x"0048", x"008C", x"00E8", x"0147", x"01A0", x"01E6", x"0211", x"0210", x"0203", x"01F3", x"01DE", x"01E7", x"01EC", x"01E0", x"01C6", x"018E", x"014B", x"0113", x"0109", x"011B", x"0126", x"0142", x"013D", x"011E", x"00F5", x"00DC", x"00A8", x"006B", x"0044", x"0011", x"FFD8", x"FFAB", x"FF76", x"FF1E", x"FED1", x"FE89", x"FE5C", x"FE3E", x"FE4F", x"FE6B", x"FE88", x"FEB2", x"FECE", x"FECE", x"FED8", x"FEC2", x"FEC0", x"FEBB", x"FEDA", x"FEF9", x"FF12", x"FF23", x"FF0B", x"FEDF", x"FEAF", x"FE7B", x"FE59", x"FE44", x"FE29", x"FDF7", x"FDB2", x"FD59", x"FCF2", x"FCB5", x"FCAB", x"FCBF", x"FCEF", x"FD38", x"FD67", x"FD94", x"FDD0", x"FE1F", x"FE54", x"FE9E", x"FED8", x"FEF7", x"FEFB", x"FEFC", x"FECE", x"FE81", x"FE2F", x"FDD8", x"FD7C", x"FD43", x"FD1C", x"FD02", x"FD00", x"FD11", x"FD23", x"FD3B", x"FD65", x"FD8A", x"FDBC", x"FE05", x"FE62", x"FEC2", x"FF2A", x"FF7C", x"FFA3", x"FFB1", x"FFA5", x"FF89", x"FF6B", x"FF4D", x"FF19", x"FEC8", x"FE60", x"FDCF", x"FD36", x"FCC6", x"FC7D", x"FC54", x"FC54", x"FC62", x"FC59", x"FC60", x"FC84", x"FCAA", x"FCC8", x"FCFB", x"FD1A", x"FD28", x"FD3C", x"FD52", x"FD4B", x"FD40", x"FD3A", x"FD34", x"FD36", x"FD53", x"FD77", x"FD96", x"FDBE", x"FDE4", x"FDF1", x"FE02", x"FE0F", x"FE15", x"FE2F", x"FE69", x"FEB6", x"FF16", x"FF71", x"FFB3", x"FFCC", x"FFC5", x"FFAD", x"FF86", x"FF74", x"FF5E", x"FF47", x"FF2C", x"FF03", x"FEC4", x"FE88", x"FE81", x"FE8A", x"FEB4", x"FEF8", x"FF27", x"FF37", x"FF53", x"FF70", x"FF7F", x"FF7D", x"FF85", x"FF60", x"FF33", x"FF04", x"FEC8", x"FE68", x"FE05", x"FD9E", x"FD2F", x"FCDB", x"FCAA", x"FC8D", x"FC86", x"FC9A", x"FCA9", x"FCAC", x"FCA8", x"FC9B", x"FC79", x"FC73", x"FC7A", x"FC92", x"FCBD", x"FCEE", x"FD01", x"FD0E", x"FD0B", x"FD05", x"FD0B", x"FD2D", x"FD4D", x"FD60", x"FD63", x"FD3D", x"FCEA", x"FCAB", x"FC88", x"FC71", x"FC7A", x"FC7E", x"FC5B", x"FC18", x"FBE4", x"FBB8", x"FB8E", x"FB7D", x"FB8C", x"FB86", x"FBA3", x"FBDF", x"FC0B", x"FC3F", x"FC74", x"FCA1", x"FCCB", x"FD00", x"FD40", x"FD72", x"FDAB", x"FDD3", x"FDDF", x"FDD3", x"FDB5", x"FD81", x"FD44", x"FD21", x"FD0B", x"FD02", x"FD16", x"FD19", x"FD0B", x"FCEE", x"FCC9", x"FCA3", x"FC92", x"FCA0", x"FCA2", x"FCA8", x"FC98", x"FC6F", x"FC2F", x"FC1B", x"FC21", x"FC4B", x"FC99", x"FCE7", x"FD07", x"FD1E", x"FD3B", x"FD47", x"FD5B", x"FD7C", x"FD8C", x"FD8D", x"FD95", x"FD9C", x"FD8B", x"FD7B", x"FD67", x"FD3A", x"FD17", x"FD02", x"FCF5", x"FCF6", x"FD06", x"FD17", x"FD15", x"FD18", x"FD1E", x"FD0F", x"FD21", x"FD37", x"FD5E", x"FD89", x"FDC4", x"FDF3", x"FE0A", x"FE28", x"FE37", x"FE4A", x"FE72", x"FEA5", x"FEC6", x"FEEC", x"FEEB", x"FEC7", x"FE93", x"FE77", x"FE5F", x"FE6B", x"FE91", x"FEA5", x"FE9F", x"FE9F", x"FEA2", x"FE9C", x"FE99", x"FEA7", x"FE80", x"FE63", x"FE39", x"FE11", x"FDCC", x"FD9A", x"FD57", x"FD0E", x"FCDC", x"FCC2", x"FCB8", x"FCC3", x"FCE8", x"FD0E", x"FD2B", x"FD56", x"FD70", x"FD7E", x"FD93", x"FDB4", x"FDDA", x"FE0D", x"FE3D", x"FE4C", x"FE3A", x"FE0E", x"FDD4", x"FDA1", x"FD82", x"FD76", x"FD6E", x"FD7A", x"FD68", x"FD4E", x"FD42", x"FD52", x"FD75", x"FDD1", x"FE34", x"FE79", x"FEA3", x"FEBC", x"FECB", x"FEBA", x"FEC2", x"FEAA", x"FE72", x"FE26", x"FDE0", x"FD7A", x"FD11", x"FCB2", x"FC4B", x"FBEE", x"FBB7", x"FBA3", x"FBAD", x"FBDD", x"FC41", x"FC9E", x"FD14", x"FD83", x"FDE4", x"FE2B", x"FE82", x"FECF", x"FF37", x"FF9F", x"000A", x"004E", x"007E", x"0091", x"0092", x"00A2", x"00B2", x"00C2", x"00C6", x"00C8", x"008E", x"004E", x"0016", x"FFF8", x"FFF2", x"001C", x"003E", x"003C", x"001A", x"0011", x"FFE3", x"FFC6", x"FFB3", x"FF8D", x"FF50", x"FF22", x"FF0F", x"FEE5", x"FED4", x"FEB7", x"FE99", x"FE69", x"FE64", x"FE5C", x"FE65", x"FE81", x"FEA2", x"FEB9", x"FED3", x"FEED", x"FEF3", x"FF03", x"FF1B", x"FF3E", x"FF6E", x"FF9F", x"FFC2", x"FFC0", x"FFAE", x"FF89", x"FF61", x"FF4A", x"FF3C", x"FF1E", x"FF0F", x"FEE4", x"FE98", x"FE4C", x"FE1D", x"FE05", x"FE1D", x"FE66", x"FEAF", x"FEDA", x"FF17", x"FF50", x"FF85", x"FFBD", x"0002", x"0016", x"0025", x"0028", x"0036", x"0015", x"0008", x"FFD4", x"FF8E", x"FF3D", x"FEFE", x"FEB4", x"FE8A", x"FE74", x"FE5F", x"FE5C", x"FE66", x"FE77", x"FE8B", x"FEB7", x"FEF0", x"FF35", x"FF8F", x"FFF5", x"004B", x"0092", x"00CB", x"00E6", x"00F7", x"0107", x"010F", x"0102", x"00F5", x"00BE", x"0050", x"FFEB", x"FF87", x"FF3C", x"FF21", x"FF38", x"FF38", x"FF3D", x"FF4E", x"FF6B", x"FF86", x"FFC5", x"FFFA", x"001A", x"0025", x"0040", x"0040", x"0042", x"0043", x"003E", x"0024", x"0021", x"0022", x"0020", x"002B", x"0045", x"004C", x"0062", x"0085", x"00A4", x"00CB", x"0108", x"0158", x"01B9", x"022D", x"02A6", x"02F4", x"0329", x"0330", x"031F", x"0306", x"02EF", x"02DB", x"02BF", x"02A4", x"0264", x"0213", x"01D7", x"01A7", x"019E", x"01C9", x"020A", x"0226", x"0241", x"0258", x"0262", x"0272", x"029C", x"02AB", x"02A1", x"0295", x"0283", x"025E", x"0236", x"020D", x"01C2", x"016D", x"012B", x"00E5", x"00B4", x"00A0", x"00A1", x"009F", x"00B5", x"00CC", x"00D7", x"00D5", x"00E8", x"00E9", x"0103", x"0129", x"014C", x"0167", x"017A", x"0188", x"0195", x"01B7", x"01DF", x"01FF", x"021F", x"021E", x"01F0", x"01A8", x"016F", x"012F", x"0115", x"011D", x"0119", x"00E5", x"00BC", x"0096", x"0074", x"0076", x"00A3", x"00B5", x"00C8", x"00F2", x"0125", x"0155", x"0199", x"01DB", x"01F7", x"0218", x"0242", x"025B", x"0279", x"029D", x"02A9", x"02A8", x"02A1", x"0298", x"0276", x"0266", x"0251", x"024B", x"024A", x"0264", x"0266", x"0262", x"024D", x"0228", x"0209", x"01F4", x"01F3", x"01E9", x"01FD", x"01E2", x"01B1", x"017B", x"0152", x"0138", x"0159", x"019F", x"01DE", x"01FB", x"022F", x"0249", x"0266", x"029A", x"02D1", x"02E2", x"02ED", x"02FB", x"02FC", x"02F6", x"0303", x"02EE", x"02C7", x"029E", x"026D", x"0234", x"020E", x"01F5", x"01CC", x"01B9", x"01AD", x"01A4", x"019F", x"01B2", x"01C6", x"01DF", x"0218", x"0254", x"028D", x"02D0", x"0301", x"0329", x"034B", x"0384", x"03AC", x"03E0", x"0413", x"040F", x"03E6", x"03B4", x"0376", x"033C", x"033B", x"0345", x"0335", x"030F", x"0300", x"02CB", x"02B9", x"02C0", x"02C4", x"02AD", x"0297", x"0281", x"0250", x"022E", x"020F", x"01E3", x"01B0", x"019A", x"0185", x"0187", x"01A5", x"01CF", x"01EB", x"021A", x"0241", x"0262", x"027D", x"02AE", x"02D0", x"0305", x"0340", x"037B", x"0394", x"039B", x"0379", x"033F", x"030D", x"02E3", x"02C1", x"02B5", x"02B0", x"0288", x"0267", x"0249", x"0236", x"0251", x"029E", x"02F7", x"0322", x"034C", x"0357", x"0349", x"034F", x"0366", x"0360", x"033A", x"031E", x"02E5", x"02A2", x"026E", x"0239", x"01EE", x"01B2", x"0186", x"0167", x"015D", x"017E", x"019D", x"01C7", x"0204", x"023B", x"0263", x"0299", x"02C1", x"02EC", x"0319", x"035F", x"0395", x"03CB", x"03FA", x"0411", x"0424", x"043C", x"0451", x"045F", x"047A", x"0479", x"044A", x"0417", x"03DC", x"03A1", x"0399", x"03C0", x"03CF", x"03B8", x"039F", x"036E", x"032D", x"0320", x"031D", x"02FD", x"02D9", x"02C5", x"02A1", x"0280", x"027D", x"026A", x"024C", x"023A", x"0233", x"0223", x"0227", x"0235", x"0235", x"0232", x"0240", x"0239", x"0238", x"0250", x"025D", x"0275", x"0297", x"02C1", x"02CE", x"02E6", x"02DC", x"02BC", x"028D", x"0266", x"0235", x"0214", x"020E", x"01E5", x"01AC", x"0174", x"0138", x"0111", x"012A", x"016E", x"0198", x"01BC", x"01DD", x"01E3", x"01EF", x"0228", x"0256", x"0270", x"0283", x"0291", x"0275", x"025F", x"0242", x"020C", x"01CF", x"018B", x"0140", x"00E8", x"00B6", x"007D", x"0055", x"004C", x"004E", x"0052", x"0079", x"00B2", x"00E6", x"0128", x"0182", x"01D2", x"021D", x"0278", x"02A8", x"02BE", x"02CC", x"02D4", x"02C2", x"02CC", x"02C2", x"0288", x"0229", x"01B6", x"012C", x"00BB", x"008C", x"007A", x"0052", x"0048", x"0031", x"001A", x"0020", x"005B", x"0085", x"00A6", x"00C9", x"00D0", x"00BD", x"00B8", x"00AF", x"009A", x"008A", x"008B", x"007E", x"008C", x"00AC", x"00CA", x"00EB", x"0123", x"0153", x"0186", x"01D8", x"022A", x"027D", x"02DE", x"034B", x"039A", x"03DF", x"0401", x"03F0", x"03B8", x"037C", x"0338", x"02FF", x"02E1", x"02C3", x"0287", x"024E", x"020A", x"01CA", x"01B7", x"01F4", x"0221", x"024F", x"0270", x"026F", x"0251", x"0262", x"0277", x"027A", x"026B", x"0262", x"022C", x"01F4", x"01C2", x"0184", x"0123", x"00D7", x"0086", x"0039", x"0003", x"FFE4", x"FFBA", x"FF9F", x"FF97", x"FF86", x"FF82", x"FF97", x"FFA1", x"FFAE", x"FFCF", x"FFF1", x"0008", x"0031", x"0050", x"005B", x"006A", x"0082", x"0089", x"00A5", x"00DA", x"00DE", x"00D3", x"009D", x"0048", x"FFD0", x"FFA6", x"FF98", x"FF7E", x"FF5F", x"FF3A", x"FEE9", x"FEA4", x"FEAB", x"FEBD", x"FECA", x"FEE7", x"FF0C", x"FF11", x"FF25", x"FF4C", x"FF55", x"FF5A", x"FF6F", x"FF82", x"FF87", x"FFA0", x"FFA4", x"FF97", x"FF8D", x"FF7B", x"FF5E", x"FF46", x"FF45", x"FF35", x"FF37", x"FF4E", x"FF5B", x"FF6F", x"FF91", x"FF9E", x"FF8F", x"FF86", x"FF72", x"FF4B", x"FF4E", x"FF5F", x"FF4F", x"FF2F", x"FEFD", x"FEA0", x"FE5C", x"FE67", x"FE93", x"FEB8", x"FEE6", x"FF00", x"FEED", x"FEF4", x"FF2F", x"FF5D", x"FF84", x"FFBA", x"FFD7", x"FFDB", x"FFEE", x"FFFB", x"FFF5", x"FFE8", x"FFE1", x"FFB3", x"FF84", x"FF51", x"FF06", x"FED0", x"FEA3", x"FE85", x"FE5F", x"FE6C", x"FE79", x"FE8E", x"FEC9", x"FF09", x"FF4B", x"FF9C", x"0002", x"004B", x"0083", x"00C6", x"00E3", x"00FF", x"0130", x"0157", x"0140", x"011E", x"00C8", x"0042", x"FFE6", x"FFBE", x"FFAD", x"FF99", x"FF9B", x"FF7B", x"FF45", x"FF3D", x"FF52", x"FF4D", x"FF4A", x"FF4A", x"FF28", x"FEFA", x"FEEA", x"FEC5", x"FE95", x"FE76", x"FE52", x"FE2B", x"FE15", x"FE08", x"FDEB", x"FDDD", x"FDD8", x"FDC6", x"FDC3", x"FDDC", x"FDFA", x"FE1A", x"FE5A", x"FE95", x"FEBE", x"FEF1", x"FF0D", x"FF00", x"FEE1", x"FEBC", x"FE7D", x"FE5A", x"FE5D", x"FE5B", x"FE4B", x"FE44", x"FE0C", x"FDC7", x"FDBF", x"FDDE", x"FE01", x"FE2F", x"FE53", x"FE38", x"FE19", x"FE20", x"FE2F", x"FE27", x"FE27", x"FE26", x"FDEF", x"FDD2", x"FDBB", x"FD8E", x"FD62", x"FD47", x"FD32", x"FD1C", x"FD1E", x"FD20", x"FD0D", x"FD0F", x"FD15", x"FD1A", x"FD36", x"FD5F", x"FD7E", x"FDAE", x"FDE3", x"FE14", x"FE40", x"FE81", x"FEAB", x"FED1", x"FEF7", x"FF16", x"FF20", x"FF53", x"FF92", x"FFB2", x"FFD1", x"FFC7", x"FF7A", x"FF22", x"FF06", x"FEFE", x"FEEE", x"FEF0", x"FEC9", x"FE63", x"FE0F", x"FDFA", x"FDDD", x"FDC4", x"FDCB", x"FDB8", x"FD86", x"FD78", x"FD71", x"FD50", x"FD3C", x"FD3E", x"FD38", x"FD3E", x"FD51", x"FD5A", x"FD4E", x"FD4B", x"FD46", x"FD2D", x"FD36", x"FD32", x"FD34", x"FD4B", x"FD68", x"FD77", x"FD94", x"FDAD", x"FDB2", x"FDAA", x"FDA4", x"FD82", x"FD57", x"FD5D", x"FD60", x"FD53", x"FD5E", x"FD3E", x"FD04", x"FCE1", x"FCF6", x"FD14", x"FD2B", x"FD5A", x"FD4A", x"FD21", x"FD20", x"FD48", x"FD64", x"FD90", x"FDC7", x"FDD3", x"FDD4", x"FDE5", x"FDE4", x"FDC9", x"FDB6", x"FD94", x"FD61", x"FD29", x"FCF2", x"FCA8", x"FC67", x"FC35", x"FC04", x"FBEC", x"FBF5", x"FC00", x"FC26", x"FC5A", x"FC8F", x"FCB1", x"FCF1", x"FD21", x"FD4B", x"FD7D", x"FDAE", x"FDC1", x"FDE1", x"FE11", x"FE2B", x"FE28", x"FE1D", x"FDCF", x"FD56", x"FD03", x"FCCE", x"FCA6", x"FC97", x"FC9E", x"FC6E", x"FC44", x"FC49", x"FC61", x"FC71", x"FC9C", x"FCB1", x"FCA6", x"FC90", x"FC95", x"FC7B", x"FC5F", x"FC55", x"FC53", x"FC52", x"FC75", x"FC94", x"FCB3", x"FCD1", x"FD01", x"FD24", x"FD6D", x"FDB8", x"FE12", x"FE66", x"FED0", x"FF19", x"FF6C", x"FFB0", x"FFE0", x"FFE7", x"FFE4", x"FFC0", x"FF82", x"FF5D", x"FF45", x"FF2B", x"FF17", x"FEFE", x"FEBB", x"FE6D", x"FE59", x"FE5A", x"FE73", x"FEA7", x"FECB", x"FEB2", x"FEA1", x"FEAF", x"FEB6", x"FEC1", x"FECC", x"FEC0", x"FE86", x"FE5C", x"FE35", x"FDF4", x"FDBD", x"FD93", x"FD73", x"FD4B", x"FD46", x"FD22", x"FCF7", x"FCCE", x"FC9E", x"FC7D", x"FC67", x"FC63", x"FC66", x"FC84", x"FCA8", x"FCD1", x"FCFD", x"FD31", x"FD4E", x"FD76", x"FDA1", x"FDBB", x"FDD5", x"FE02", x"FE2F", x"FE4C", x"FE67", x"FE5F", x"FE15", x"FDCE", x"FDB0", x"FD93", x"FD95", x"FDA9", x"FDA3", x"FD64", x"FD5E", x"FD68", x"FD7E", x"FDA3", x"FDD4", x"FDE6", x"FDD9", x"FDF7", x"FDFF", x"FDF7", x"FDF3", x"FDF9", x"FDFE", x"FE11", x"FE3B", x"FE54", x"FE62", x"FE6E", x"FE68", x"FE61", x"FE64", x"FE67", x"FE73", x"FE8E", x"FEB2", x"FECB", x"FEEB", x"FF06", x"FF05", x"FF05", x"FEF4", x"FECE", x"FEA0", x"FE89", x"FE5B", x"FE37", x"FE10", x"FDD6", x"FD84", x"FD56", x"FD4B", x"FD4E", x"FD76", x"FDA6", x"FDB7", x"FDB8", x"FDE3", x"FE17", x"FE58", x"FEB0", x"FF06", x"FF32", x"FF5F", x"FF84", x"FF97", x"FF8D", x"FF90", x"FF7C", x"FF61", x"FF46", x"FF1E", x"FEE1", x"FE99", x"FE59", x"FE19", x"FDF7", x"FDF7", x"FE05", x"FE2E", x"FE6C", x"FEAC", x"FEEF", x"FF52", x"FFAB", x"0009", x"0068", x"00B2", x"00E9", x"0118", x"0143", x"0157", x"0153", x"0140", x"00F6", x"0097", x"004D", x"0011", x"FFEA", x"FFE3", x"FFE1", x"FFB2", x"FF95", x"FF85", x"FF82", x"FF80", x"FFA2", x"FF9F", x"FF8A", x"FF77", x"FF74", x"FF51", x"FF3C", x"FF2C", x"FF10", x"FF02", x"FF08", x"FF16", x"FF0E", x"FF14", x"FF14", x"FF15", x"FF2F", x"FF5D", x"FF8F", x"FFC3", x"0000", x"002B", x"0056", x"007E", x"009E", x"00A4", x"00A7", x"0094", x"0078", x"0064", x"0058", x"0049", x"0043", x"0037", x"000F", x"FFEE", x"FFDD", x"FFD6", x"FFE3", x"0002", x"0009", x"FFF8", x"FFEE", x"0001", x"0009", x"0032", x"0060", x"0070", x"006A", x"0079", x"0084", x"007B", x"0078", x"007B", x"005E", x"0058", x"0055", x"0050", x"0037", x"0026", x"0013", x"FFFE", x"0007", x"001D", x"0036", x"0066", x"0092", x"00C7", x"00F6", x"0134", x"0163", x"019D", x"01DF", x"0211", x"024E", x"0288", x"02BE", x"02E4", x"0308", x"0302", x"02C9", x"028C", x"0249", x"020C", x"01E3", x"01D8", x"01A0", x"0157", x"0130", x"010B", x"00FD", x"010D", x"0130", x"0126", x"012B", x"0139", x"0140", x"012F", x"0139", x"013A", x"0133", x"0153", x"0175", x"0186", x"0184", x"0179", x"0155", x"0132", x"0121", x"0113", x"010B", x"0110", x"0120", x"012A", x"0149", x"0165", x"0178", x"018C", x"019B", x"019D", x"01A0", x"01AC", x"01A7", x"01A6", x"01A1", x"0183", x"0157", x"0134", x"011B", x"0107", x"0112", x"011A", x"0101", x"00ED", x"00E7", x"00F1", x"010C", x"014D", x"0183", x"01A5", x"01CD", x"01EE", x"01F6", x"01F3", x"01F3", x"01DB", x"01C4", x"01B6", x"01A3", x"0173", x"014E", x"0112", x"00DA", x"00B6", x"00AC", x"00AB", x"00C5", x"00EB", x"0111", x"0136", x"0175", x"01A7", x"01E1", x"021E", x"0255", x"027F", x"02A5", x"02C2", x"02CB", x"02C3", x"02AD", x"026E", x"0225", x"01E5", x"01A5", x"017A", x"0165", x"014F", x"0122", x"0111", x"0108", x"010B", x"0120", x"0148", x"0151", x"0147", x"0149", x"013A", x"0121", x"0111", x"0109", x"00F7", x"010D", x"013C", x"0178", x"01B0", x"01FB", x"0229", x"0253", x"028D", x"02CD", x"030E", x"0356", x"039E", x"03CF", x"03FD", x"042D", x"044C", x"045A", x"0467", x"0455", x"0440", x"0424", x"0419", x"0402", x"03F7", x"03E3", x"03B8", x"0397", x"0375", x"0368", x"0364", x"037F", x"037A", x"0367", x"035B", x"033C", x"0325", x"0310", x"0306", x"02D5", x"02AA", x"0286", x"024F", x"0223", x"01F8", x"01DF", x"01B8", x"01B3", x"01B9", x"01A9", x"01A8", x"0190", x"0175", x"0151", x"0148", x"013D", x"013F", x"0148", x"015B", x"0159", x"0177", x"018C", x"01B0", x"01DA", x"020B", x"0233", x"025C", x"028F", x"02BA", x"02DD", x"0308", x"02FD", x"02DF", x"02B4", x"0278", x"0247", x"0228", x"0223", x"01FA", x"01DE", x"01CA", x"01B4", x"01B2", x"01CC", x"01E8", x"01E4", x"01EE", x"01FB", x"01E2", x"01DB", x"01C9", x"01BC", x"01A7", x"01BF", x"01DC", x"01F3", x"0214", x"0220", x"0218", x"020F", x"0210", x"0211", x"0221", x"023E", x"0253", x"0267", x"0281", x"0291", x"029E", x"029C", x"02A0", x"0284", x"0280", x"0272", x"0264", x"0258", x"0243", x"0214", x"01DA", x"01A4", x"0164", x"0139", x"0129", x"011A", x"010D", x"010E", x"0127", x"0149", x"018A", x"01E6", x"0230", x"0272", x"02B5", x"02E3", x"02FC", x"030E", x"0312", x"0301", x"02F2", x"02E0", x"02C7", x"02A3", x"0285", x"0255", x"0224", x"020A", x"01FE", x"020B", x"022F", x"0268", x"0296", x"02D0", x"0318", x"035C", x"03A5", x"03F2", x"0424", x"0449", x"0464", x"0471", x"046A", x"0460", x"0438", x"03FA", x"03A9", x"035B", x"030C", x"02D6", x"02BD", x"029D", x"0284", x"0272", x"025F", x"0250", x"0255", x"0262", x"025B", x"0253", x"0241", x"0216", x"01DE", x"01A1", x"0162", x"0117", x"00F4", x"00D1", x"00CE", x"00CA", x"00E6", x"00DD", x"00E9", x"00F6", x"010B", x"012B", x"0160", x"0191", x"01B1", x"01DF", x"020A", x"0234", x"0259", x"0279", x"027D", x"0272", x"0268", x"0264", x"024D", x"0249", x"022F", x"0206", x"01DD", x"01B3", x"018A", x"0173", x"0161", x"0150", x"013F", x"012F", x"0128", x"0120", x"0138", x"0151", x"0170", x"018F", x"01B0", x"01BA", x"01C5", x"01BF", x"01B8", x"019E", x"019A", x"0186", x"0172", x"0166", x"014A", x"0123", x"00FD", x"00E1", x"00C4", x"00C1", x"00C7", x"00CB", x"00CD", x"00E4", x"0102", x"0126", x"0162", x"019E", x"01D2", x"020D", x"024E", x"0280", x"02AB", x"02C8", x"02C3", x"02A3", x"027B", x"0242", x"0211", x"01F2", x"01DA", x"01B7", x"0191", x"016F", x"013A", x"011B", x"0109", x"00F9", x"00E8", x"00E6", x"00E3", x"00D7", x"00D4", x"00CC", x"00BD", x"00B3", x"00BC", x"00C8", x"00D3", x"00E9", x"00E6", x"00CC", x"00B9", x"009C", x"007A", x"0075", x"0068", x"0063", x"0062", x"007C", x"00A5", x"00CB", x"0106", x"012B", x"014C", x"0163", x"018A", x"0196", x"01AA", x"019D", x"0182", x"0146", x"0109", x"00C0", x"0089", x"005D", x"0039", x"0010", x"FFF6", x"FFDC", x"FFD1", x"FFE7", x"0013", x"0045", x"0085", x"00C2", x"00EB", x"010C", x"0112", x"010C", x"00E8", x"00C7", x"00A2", x"0074", x"0048", x"0019", x"FFD6", x"FF8A", x"FF4A", x"FF0D", x"FEDE", x"FED0", x"FEC7", x"FEBC", x"FEC5", x"FEDC", x"FEFF", x"FF29", x"FF64", x"FF8E", x"FFB4", x"FFDC", x"0008", x"0024", x"0044", x"0045", x"0030", x"FFFD", x"FFBC", x"FF7B", x"FF3B", x"FF16", x"FEED", x"FED0", x"FEB8", x"FE9B", x"FE89", x"FE86", x"FE89", x"FE8A", x"FE91", x"FE93", x"FE86", x"FE75", x"FE67", x"FE43", x"FE34", x"FE2F", x"FE4B", x"FE6E", x"FEB8", x"FF02", x"FF3E", x"FF7D", x"FFB6", x"FFE4", x"0014", x"004F", x"007B", x"008D", x"00B2", x"00CB", x"00E0", x"00F6", x"0109", x"0101", x"00F4", x"00ED", x"00F2", x"00E7", x"00EB", x"00D9", x"00BE", x"0091", x"007C", x"0051", x"0045", x"0036", x"001F", x"0005", x"FFDB", x"FFB3", x"FF88", x"FF6D", x"FF5E", x"FF4F", x"FF4C", x"FF47", x"FF2C", x"FF13", x"FEE9", x"FEBC", x"FE8F", x"FE76", x"FE61", x"FE56", x"FE5A", x"FE55", x"FE41", x"FE32", x"FE19", x"FDF6", x"FDDE", x"FDC9", x"FDA8", x"FD92", x"FD8F", x"FD9A", x"FDB0", x"FDE0", x"FE08", x"FE26", x"FE4F", x"FE84", x"FEB7", x"FEF2", x"FF27", x"FF3B", x"FF32", x"FF1D", x"FEF2", x"FECD", x"FEB3", x"FEA1", x"FE85", x"FE71", x"FE5B", x"FE3A", x"FE35", x"FE34", x"FE3B", x"FE3C", x"FE4F", x"FE50", x"FE50", x"FE46", x"FE38", x"FE17", x"FE07", x"FE0B", x"FE17", x"FE3A", x"FE62", x"FE7D", x"FE86", x"FE93", x"FE92", x"FE88", x"FE96", x"FE8F", x"FE88", x"FE7A", x"FE79", x"FE6F", x"FE73", x"FE7A", x"FE73", x"FE62", x"FE55", x"FE4F", x"FE3E", x"FE3B", x"FE26", x"FDF9", x"FDBB", x"FD7A", x"FD39", x"FD0B", x"FCFB", x"FCF9", x"FCF3", x"FD08", x"FD0E", x"FD29", x"FD50", x"FD93", x"FDD0", x"FE1C", x"FE6B", x"FEAC", x"FED9", x"FEFE", x"FEF6", x"FEDF", x"FEB9", x"FE98", x"FE6F", x"FE52", x"FE34", x"FE05", x"FDDF", x"FDB6", x"FD8D", x"FD76", x"FD7D", x"FD82", x"FDA0", x"FDCA", x"FE04", x"FE40", x"FE8F", x"FEDC", x"FF0D", x"FF2E", x"FF4A", x"FF56", x"FF58", x"FF60", x"FF4B", x"FF1C", x"FEE1", x"FE9B", x"FE5C", x"FE2F", x"FE22", x"FE0E", x"FE01", x"FDF4", x"FDD6", x"FDBF", x"FDBE", x"FDB1", x"FDB3", x"FDAB", x"FDA6", x"FD89", x"FD66", x"FD3D", x"FD01", x"FCD0", x"FCB5", x"FCA7", x"FCB0", x"FCD4", x"FCF3", x"FD11", x"FD2F", x"FD47", x"FD4D", x"FD6A", x"FD88", x"FD9C", x"FDBE", x"FDDC", x"FDFF", x"FE12", x"FE40", x"FE53", x"FE53", x"FE50", x"FE55", x"FE50", x"FE5E", x"FE72", x"FE67", x"FE46", x"FE20", x"FDED", x"FDC6", x"FDB0", x"FDAB", x"FD9E", x"FD93", x"FD88", x"FD77", x"FD6F", x"FD80", x"FD9D", x"FDC5", x"FE01", x"FE3D", x"FE61", x"FE81", x"FE7E", x"FE68", x"FE4C", x"FE2D", x"FE17", x"FE03", x"FDFD", x"FDE8", x"FDDD", x"FDC5", x"FDA6", x"FD83", x"FD74", x"FD62", x"FD5D", x"FD64", x"FD79", x"FD88", x"FDBD", x"FDFE", x"FE3B", x"FE75", x"FEB0", x"FED9", x"FEFA", x"FF20", x"FF3E", x"FF30", x"FF17", x"FEEF", x"FEB4", x"FE8F", x"FE7A", x"FE69", x"FE4A", x"FE37", x"FE0C", x"FDE2", x"FDCC", x"FDCA", x"FDCF", x"FDE9", x"FE10", x"FE38", x"FE50", x"FE73", x"FE71", x"FE6B", x"FE65", x"FE6D", x"FE73", x"FE97", x"FEAF", x"FEC6", x"FECF", x"FEC9", x"FEAB", x"FE86", x"FE63", x"FE3E", x"FE20", x"FE19", x"FE16", x"FE1D", x"FE47", x"FE77", x"FE9F", x"FED3", x"FEF9", x"FF1C", x"FF31", x"FF61", x"FF62", x"FF51", x"FF26", x"FEE1", x"FE8E", x"FE4D", x"FE1C", x"FDEF", x"FDC4", x"FDA9", x"FD7F", x"FD6C", x"FD75", x"FD99", x"FDCB", x"FE1A", x"FE6C", x"FEB3", x"FEDE", x"FF00", x"FEEC", x"FED6", x"FEA4", x"FE81", x"FE4F", x"FE34", x"FE11", x"FE01", x"FDEE", x"FDDF", x"FDC4", x"FDB8", x"FDA0", x"FD93", x"FD92", x"FD9E", x"FDA4", x"FDBD", x"FDF0", x"FE19", x"FE4D", x"FE7F", x"FEAF", x"FEC8", x"FEFB", x"FF1C", x"FF2A", x"FF1D", x"FEFE", x"FEBE", x"FE88", x"FE62", x"FE51", x"FE42", x"FE3E", x"FE36", x"FE19", x"FE06", x"FE00", x"FDFB", x"FE0C", x"FE2A", x"FE4C", x"FE60", x"FE6D", x"FE69", x"FE4F", x"FE3E", x"FE35", x"FE42", x"FE6C", x"FEA8", x"FEF0", x"FF39", x"FF81", x"FFB3", x"FFD6", x"0000", x"0014", x"002E", x"0047", x"0062", x"006D", x"008C", x"00AF", x"00C8", x"00E3", x"00F6", x"0103", x"0102", x"0114", x"0120", x"010E", x"00FD", x"00D9", x"00AE", x"0087", x"0077", x"005E", x"0047", x"001F", x"FFF1", x"FFB0", x"FF7A", x"FF57", x"FF3C", x"FF45", x"FF59", x"FF75", x"FF8D", x"FF95", x"FF8D", x"FF72", x"FF61", x"FF4F", x"FF54", x"FF5F", x"FF71", x"FF7E", x"FF87", x"FF83", x"FF6D", x"FF53", x"FF38", x"FF17", x"FF05", x"FEFE", x"FEF9", x"FEFC", x"FF1D", x"FF49", x"FF7E", x"FFC5", x"0006", x"0036", x"006D", x"00A9", x"00CE", x"00E3", x"00ED", x"00CE", x"00AB", x"0088", x"007C", x"0061", x"0051", x"0031", x"FFFA", x"FFC3", x"FFA0", x"FF85", x"FF82", x"FF8A", x"FFA7", x"FFAF", x"FFC8", x"FFC9", x"FFC3", x"FFB0", x"FFAA", x"FFA4", x"FFB4", x"FFC7", x"FFE8", x"FFFD", x"001C", x"002D", x"003B", x"0045", x"0041", x"003A", x"0034", x"002B", x"0025", x"0026", x"0042", x"005B", x"0082", x"00AE", x"00BB", x"00BB", x"00BA", x"00AB", x"0097", x"0077", x"0054", x"0016", x"FFDE", x"FFC6", x"FFB7", x"FFBE", x"FFD4", x"FFE4", x"FFE6", x"FFF0", x"000D", x"0038", x"0077", x"00D8", x"0135", x"0195", x"01E6", x"0221", x"0232", x"0229", x"0218", x"01F6", x"01E2", x"01CD", x"01C1", x"01B7", x"01AB", x"01A0", x"0191", x"0185", x"0175", x"0179", x"0188", x"019C", x"01BE", x"01EB", x"0215", x"0249", x"027D", x"02B4", x"02C8", x"02DA", x"02E4", x"02E5", x"02D6", x"02CE", x"02AB", x"0271", x"024A", x"0228", x"021A", x"020F", x"0219", x"0204", x"01E4", x"01C8", x"01A9", x"0190", x"0181", x"0178", x"016D", x"014E", x"0136", x"00FA", x"00B8", x"0075", x"0040", x"0022", x"0022", x"0038", x"0060", x"008F", x"00C6", x"00F6", x"012C", x"0155", x"017E", x"01A3", x"01C3", x"01DD", x"01E9", x"0203", x"0210", x"022F", x"0255", x"0282", x"029B", x"02BF", x"02E2", x"02F0", x"02FD", x"02FE", x"02DE", x"02AE", x"028A", x"026C", x"0256", x"024B", x"023A", x"0211", x"01E0", x"01BC", x"01A6", x"01A9", x"01D0", x"020C", x"024C", x"028B", x"02BB", x"02C3", x"02B7", x"0299", x"0278", x"025B", x"024D", x"023B", x"0232", x"0224", x"0216", x"0202", x"01F3", x"01D9", x"01BD", x"01B0", x"0198", x"018F", x"018E", x"01A9", x"01CE", x"020F", x"0267", x"02A5", x"02D7", x"02FD", x"031A", x"031F", x"0336", x"0338", x"031E", x"02FF", x"02E1", x"02D3", x"02B3", x"02B3", x"0291", x"025E", x"022F", x"0209", x"01F4", x"01EC", x"0204", x"021B", x"0231", x"024C", x"0254", x"0250", x"0238", x"022E", x"0223", x"022D", x"0240", x"0258", x"0272", x"0283", x"0297", x"02A3", x"02A6", x"029E", x"0295", x"0288", x"027E", x"0271", x"0286", x"0291", x"02BB", x"02FB", x"0340", x"036C", x"0390", x"03A2", x"039B", x"038D", x"037E", x"0352", x"0305", x"02B2", x"026F", x"0227", x"0200", x"01F2", x"01DB", x"01C2", x"01BE", x"01C5", x"01E0", x"0211", x"0260", x"02A7", x"02F1", x"0337", x"035A", x"0356", x"0336", x"02F7", x"02AB", x"0262", x"0217", x"01DF", x"01AC", x"018B", x"0178", x"016C", x"0163", x"0153", x"0154", x"014B", x"0152", x"015E", x"017A", x"01A3", x"01CF", x"021F", x"0259", x"0281", x"02A4", x"02B2", x"02AB", x"02AD", x"02B0", x"0299", x"0272", x"0253", x"023C", x"0221", x"022C", x"0229", x"021A", x"01EF", x"01D3", x"01A8", x"018B", x"0185", x"0187", x"018C", x"0194", x"0198", x"0186", x"016E", x"0151", x"0143", x"014C", x"016B", x"01A0", x"01D5", x"0216", x"0247", x"027D", x"02A5", x"02C6", x"02D1", x"02E9", x"02ED", x"02F3", x"02FC", x"0311", x"031D", x"0349", x"0375", x"0396", x"039E", x"03A7", x"0397", x"0389", x"0385", x"0380", x"0367", x"033C", x"0321", x"02FA", x"02DE", x"02D1", x"02B7", x"0281", x"0247", x"0208", x"01CE", x"01A6", x"019C", x"019E", x"01B1", x"01CA", x"01DA", x"01DB", x"01C4", x"01B0", x"018D", x"017B", x"0170", x"015E", x"015A", x"014B", x"0136", x"0129", x"0118", x"00F9", x"00EA", x"00CA", x"00B9", x"0099", x"0097", x"0098", x"00B7", x"00F5", x"0147", x"018F", x"01CA", x"0200", x"0218", x"022B", x"0247", x"024C", x"023A", x"0224", x"020B", x"01EE", x"01D6", x"01CC", x"01A1", x"016A", x"0131", x"00FD", x"00DA", x"00CE", x"00E5", x"00F9", x"0118", x"013D", x"0149", x"0156", x"014A", x"0148", x"0139", x"013E", x"0139", x"0143", x"0142", x"014B", x"0143", x"0146", x"013B", x"0120", x"0106", x"00DF", x"00AF", x"008E", x"007B", x"0073", x"0090", x"00BE", x"00F2", x"0113", x"0123", x"0126", x"0104", x"00F2", x"00E2", x"00B9", x"0088", x"0058", x"0025", x"FFF6", x"FFEF", x"FFEF", x"FFEF", x"FFE8", x"FFF4", x"FFF9", x"0012", x"004B", x"0094", x"00E4", x"0137", x"0184", x"01B5", x"01CA", x"01CC", x"01B0", x"018F", x"0169", x"0149", x"0121", x"0109", x"00EB", x"00D8", x"00CD", x"00C6", x"00C3", x"00BF", x"00B9", x"00B0", x"00AF", x"00B6", x"00C6", x"00E9", x"0114", x"0140", x"0155", x"016D", x"0167", x"015D", x"015E", x"015F", x"0149", x"0131", x"0111", x"00E9", x"00D0", x"00C9", x"00CC", x"00B0", x"009F", x"0079", x"004E", x"002A", x"001D", x"000B", x"FFFB", x"FFF1", x"FFD3", x"FFAA", x"FF74", x"FF3D", x"FF01", x"FEE1", x"FED1", x"FEE1", x"FEF7", x"FF25", x"FF50", x"FF7D", x"FFAC", x"FFD4", x"FFE4", x"FFF4", x"FFE6", x"FFD0", x"FFB9", x"FFA6", x"FFA0", x"FFB3", x"FFCB", x"FFED", x"0000", x"0019", x"001A", x"0021", x"002F", x"0030", x"0020", x"000C", x"FFEE", x"FFCC", x"FFB9", x"FFB1", x"FF9D", x"FF79", x"FF4F", x"FF20", x"FEEE", x"FEE3", x"FEF0", x"FF0C", x"FF40", x"FF77", x"FF9F", x"FFB7", x"FFBC", x"FFAF", x"FF90", x"FF7A", x"FF65", x"FF51", x"FF4A", x"FF3A", x"FF2B", x"FF1D", x"FF0E", x"FEFD", x"FEE8", x"FED5", x"FEBB", x"FEA4", x"FE96", x"FE9E", x"FEB0", x"FEE9", x"FF1E", x"FF51", x"FF7C", x"FF90", x"FF92", x"FF9C", x"FFA3", x"FFAB", x"FFA2", x"FFA0", x"FF97", x"FF8B", x"FF97", x"FFAA", x"FF9F", x"FF97", x"FF76", x"FF4E", x"FF25", x"FF1C", x"FF19", x"FF21", x"FF2E", x"FF44", x"FF49", x"FF4E", x"FF51", x"FF4E", x"FF49", x"FF58", x"FF5B", x"FF6F", x"FF6F", x"FF7B", x"FF70", x"FF74", x"FF6A", x"FF65", x"FF50", x"FF34", x"FF10", x"FEEA", x"FEDA", x"FED4", x"FEF8", x"FF2B", x"FF6D", x"FFA6", x"FFD6", x"FFE0", x"FFDD", x"FFC9", x"FFB3", x"FF83", x"FF4C", x"FF0A", x"FEB7", x"FE71", x"FE45", x"FE27", x"FE04", x"FDF3", x"FDDB", x"FDC7", x"FDBF", x"FDD9", x"FE00", x"FE34", x"FE7B", x"FEB8", x"FEDF", x"FEF6", x"FEF0", x"FECA", x"FE97", x"FE62", x"FE29", x"FDFB", x"FDD9", x"FDBC", x"FDB4", x"FDB1", x"FDBC", x"FDC6", x"FDCD", x"FDD2", x"FDD0", x"FDD8", x"FDE2", x"FDF9", x"FE1E", x"FE49", x"FE6F", x"FE8E", x"FE96", x"FE8D", x"FE75", x"FE68", x"FE59", x"FE46", x"FE41", x"FE31", x"FE24", x"FE1F", x"FE36", x"FE37", x"FE3B", x"FE30", x"FE1B", x"FDF5", x"FDDE", x"FDD5", x"FDC3", x"FDC1", x"FDC0", x"FDBD", x"FDAE", x"FDAB", x"FD98", x"FD90", x"FD8C", x"FDA4", x"FDBD", x"FDE6", x"FE14", x"FE3B", x"FE62", x"FE8D", x"FEB4", x"FED8", x"FEF0", x"FF05", x"FF0B", x"FF1A", x"FF29", x"FF46", x"FF71", x"FF9A", x"FFC6", x"FFDE", x"FFF0", x"FFE6", x"FFDF", x"FFCA", x"FFB0", x"FF84", x"FF5C", x"FF24", x"FEED", x"FEC8", x"FEAB", x"FE8E", x"FE6B", x"FE47", x"FE12", x"FDDE", x"FDC1", x"FDB4", x"FDB8", x"FDDB", x"FDFE", x"FE23", x"FE33", x"FE3F", x"FE26", x"FE0E", x"FDED", x"FDCE", x"FDB3", x"FD9D", x"FD8E", x"FD7A", x"FD70", x"FD6C", x"FD66", x"FD68", x"FD60", x"FD50", x"FD39", x"FD2B", x"FD1D", x"FD31", x"FD59", x"FD96", x"FDDB", x"FE1C", x"FE53", x"FE70", x"FE93", x"FEAE", x"FEBC", x"FEC9", x"FED0", x"FEC5", x"FEBB", x"FEB1", x"FEA7", x"FE83", x"FE60", x"FE2A", x"FDEF", x"FDBD", x"FDA2", x"FD94", x"FD91", x"FDA4", x"FDB2", x"FDBD", x"FDC5", x"FDC5", x"FDC1", x"FDB9", x"FDBB", x"FDC3", x"FDCB", x"FDD5", x"FDDB", x"FDD7", x"FDD5", x"FDCE", x"FDC8", x"FDB9", x"FDA8", x"FD8C", x"FD7C", x"FD71", x"FD74", x"FD90", x"FDB5", x"FDE9", x"FE1B", x"FE40", x"FE56", x"FE53", x"FE4A", x"FE32", x"FE06", x"FDE0", x"FDA9", x"FD6D", x"FD44", x"FD29", x"FD21", x"FD1D", x"FD2B", x"FD36", x"FD49", x"FD6C", x"FDA3", x"FDE8", x"FE3A", x"FE99", x"FEEC", x"FF33", x"FF6B", x"FF84", x"FF86", x"FF76", x"FF57", x"FF3A", x"FF12", x"FEF2", x"FED0", x"FEBA", x"FEAF", x"FEB0", x"FEB7", x"FEC3", x"FEC4", x"FECA", x"FEC9", x"FED0", x"FEDD", x"FEFD", x"FF25", x"FF52", x"FF83", x"FFA1", x"FFB5", x"FFB4", x"FFB8", x"FFAC", x"FF9C", x"FF8B", x"FF6E", x"FF55", x"FF3F", x"FF39", x"FF20", x"FF0E", x"FEE5", x"FEBB", x"FE80", x"FE56", x"FE2D", x"FE0F", x"FDFF", x"FDF6", x"FDF5", x"FDE1", x"FDDD", x"FDBE", x"FDA7", x"FD9B", x"FD9A", x"FDB1", x"FDCA", x"FDF5", x"FE17", x"FE3D", x"FE5E", x"FE82", x"FE9B", x"FEB1", x"FEBA", x"FEB5", x"FEB0", x"FEB0", x"FEBB", x"FED7", x"FF05", x"FF33", x"FF61", x"FF86", x"FF9B", x"FFAB", x"FFB0", x"FFAE", x"FFA5", x"FF93", x"FF7F", x"FF66", x"FF5C", x"FF54", x"FF48", x"FF3D", x"FF28", x"FF0C", x"FEF3", x"FEDE", x"FED8", x"FEDE", x"FEF7", x"FF1C", x"FF38", x"FF5D", x"FF64", x"FF6C", x"FF62", x"FF57", x"FF4B", x"FF39", x"FF34", x"FF1A", x"FF0B", x"FEEF", x"FEDF", x"FEC8", x"FEC5", x"FEB9", x"FEB0", x"FE9F", x"FE94", x"FE86", x"FE8F", x"FEA8", x"FED3", x"FEF8", x"FF27", x"FF45", x"FF5C", x"FF70", x"FF81", x"FF8E", x"FF98", x"FFA3", x"FFB0", x"FFBB", x"FFDB", x"FFED", x"FFF7", x"FFEF", x"FFD8", x"FFAD", x"FF81", x"FF5B", x"FF3F", x"FF27", x"FF2B", x"FF2C", x"FF3A", x"FF48", x"FF5C", x"FF65", x"FF7D", x"FF93", x"FFB0", x"FFD0", x"FFEA", x"0000", x"0007", x"0011", x"0012", x"0015", x"0016", x"000C", x"FFFD", x"FFED", x"FFE1", x"FFE8", x"FFFD", x"002A", x"005F", x"009C", x"00CB", x"00F1", x"00FF", x"0100", x"00F6", x"00D7", x"00B4", x"008C", x"0058", x"0039", x"0019", x"0006", x"FFEE", x"FFDD", x"FFC4", x"FFB4", x"FFAC", x"FFBF", x"FFCF", x"0002", x"002F", x"0063", x"0085", x"0093", x"0089", x"0061", x"0035", x"0003", x"FFD1", x"FFAF", x"FF8D", x"FF77", x"FF5B", x"FF5A", x"FF52", x"FF64", x"FF79", x"FF90", x"FF9C", x"FFA9", x"FFAD", x"FFB9", x"FFC7", x"FFEC", x"000A", x"0032", x"0049", x"0058", x"0058", x"0058", x"004F", x"0048", x"0049", x"0048", x"0057", x"0068", x"0083", x"0091", x"0093", x"008C", x"0072", x"0055", x"0040", x"0028", x"0018", x"000D", x"000D", x"000A", x"000D", x"0009", x"0006", x"FFF4", x"FFFC", x"FFFF", x"0011", x"0031", x"0054", x"0075", x"0096", x"00C0", x"00E6", x"0117", x"0147", x"016B", x"017A", x"0187", x"0185", x"018D", x"01A1", x"01C5", x"01E6", x"020F", x"0231", x"023B", x"0247", x"0240", x"022E", x"0212", x"01F6", x"01D7", x"01BF", x"01BA", x"01B6", x"01B1", x"01A1", x"018D", x"0164", x"0147", x"012C", x"0120", x"011C", x"012D", x"013C", x"014A", x"0152", x"014E", x"0132", x"0111", x"00EC", x"00C3", x"00A8", x"0095", x"0086", x"007B", x"007D", x"0082", x"0095", x"00AD", x"00CE", x"00D1", x"00DC", x"00D0", x"00CC", x"00C8", x"00E1", x"00FF", x"012C", x"015D", x"018A", x"01A7", x"01C4", x"01DB", x"01E0", x"01E9", x"01EB", x"01E5", x"01E4", x"01F2", x"01EB", x"01E7", x"01D5", x"01B6", x"0192", x"0173", x"016A", x"0159", x"0161", x"016A", x"0176", x"017C", x"018E", x"0190", x"018B", x"018C", x"0189", x"018D", x"0194", x"01A1", x"0198", x"018C", x"0177", x"015E", x"0148", x"0143", x"013C", x"0134", x"0135", x"012F", x"0133", x"014A", x"016D", x"019D", x"01D1", x"0208", x"0222", x"0234", x"022E", x"0212", x"01E2", x"01AF", x"0176", x"013D", x"0123", x"0117", x"0115", x"011B", x"012B", x"012F", x"013F", x"0161", x"0187", x"01BA", x"01F7", x"023E", x"0279", x"02B7", x"02EE", x"0301", x"0308", x"0302", x"02ED", x"02DB", x"02CA", x"02B8", x"029A", x"0280", x"0267", x"0255", x"0248", x"0250", x"0248", x"0246", x"0235", x"021E", x"0210", x"0209", x"0215", x"022D", x"024B", x"026B", x"0275", x"0283", x"027E", x"026F", x"0268", x"0252", x"0248", x"0241", x"024E", x"025C", x"0264", x"025B", x"024A", x"020F", x"01E9", x"01BB", x"019A", x"017F", x"0176", x"016A", x"015C", x"015E", x"0154", x"0148", x"013C", x"0139", x"0137", x"0142", x"0159", x"0170", x"0177", x"0184", x"018A", x"0191", x"01AB", x"01C5", x"01D6", x"01E6", x"01E9", x"01EB", x"01EB", x"0209", x"0224", x"0259", x"0282", x"02AA", x"02BB", x"02C2", x"02C1", x"02A7", x"0292", x"0273", x"024C", x"0235", x"0229", x"022A", x"0222", x"0225", x"0211", x"01F4", x"01E5", x"01D7", x"01CE", x"01D1", x"01DF", x"01EB", x"01FE", x"021E", x"0238", x"0243", x"0251", x"024E", x"024B", x"023F", x"023A", x"0222", x"01FE", x"01E2", x"01BB", x"01A4", x"019C", x"0196", x"018B", x"017E", x"0166", x"0147", x"0133", x"012C", x"0131", x"0151", x"0173", x"019B", x"01BA", x"01DA", x"01F3", x"0202", x"0228", x"0235", x"0249", x"0262", x"027A", x"028C", x"0293", x"028F", x"0265", x"0238", x"020E", x"01E7", x"01C7", x"01BE", x"01B8", x"01B7", x"01C2", x"01DE", x"01E8", x"0201", x"0212", x"0224", x"0231", x"024B", x"025A", x"0267", x"0263", x"0261", x"024D", x"0247", x"0240", x"023D", x"0233", x"022B", x"021A", x"020A", x"0211", x"0212", x"022E", x"024C", x"026A", x"0279", x"0283", x"027B", x"0268", x"024C", x"0231", x"01FF", x"01D1", x"01B4", x"018D", x"017B", x"0161", x"014E", x"012B", x"0115", x"0111", x"0112", x"0122", x"0144", x"0165", x"017C", x"019D", x"01A7", x"01A0", x"0189", x"016C", x"0149", x"0129", x"0113", x"00F9", x"00DF", x"00B9", x"00A8", x"0094", x"0091", x"009E", x"00A2", x"00A7", x"00A1", x"0090", x"0082", x"006E", x"006A", x"0075", x"0085", x"00A3", x"00B2", x"00C9", x"00CB", x"00D0", x"00D8", x"00DB", x"00E3", x"00EC", x"0107", x"011A", x"0133", x"0149", x"0144", x"0133", x"011E", x"0108", x"00F2", x"00DD", x"00D7", x"00BC", x"00B1", x"00A4", x"0094", x"007D", x"006D", x"0063", x"005E", x"006D", x"0083", x"009E", x"00B1", x"00C8", x"00E2", x"00F7", x"0115", x"0136", x"0147", x"0156", x"0154", x"014C", x"0147", x"0149", x"0154", x"0170", x"0184", x"01A1", x"01A1", x"01A3", x"018F", x"0173", x"0158", x"0130", x"010E", x"00EF", x"00E6", x"00DA", x"00D8", x"00D7", x"00BE", x"00AC", x"0094", x"008B", x"0079", x"0078", x"0078", x"006F", x"0072", x"0074", x"0070", x"0060", x"0050", x"003F", x"0028", x"001F", x"0018", x"0007", x"FFF6", x"FFE9", x"FFDC", x"FFDB", x"FFDE", x"FFEC", x"FFEA", x"FFEF", x"FFE6", x"FFDF", x"FFDE", x"FFE0", x"FFF0", x"0004", x"0023", x"003F", x"0059", x"0071", x"0078", x"0081", x"0086", x"0078", x"006F", x"005F", x"004D", x"003E", x"0029", x"0014", x"FFE7", x"FFBA", x"FF93", x"FF62", x"FF45", x"FF2E", x"FF25", x"FF18", x"FF19", x"FF26", x"FF20", x"FF2A", x"FF2D", x"FF36", x"FF3D", x"FF4F", x"FF5D", x"FF5B", x"FF54", x"FF44", x"FF2A", x"FF15", x"FF05", x"FEF6", x"FEE5", x"FEDD", x"FED8", x"FEE3", x"FEF0", x"FF11", x"FF34", x"FF5C", x"FF79", x"FF90", x"FF8D", x"FF7E", x"FF58", x"FF2C", x"FEF9", x"FEC2", x"FE97", x"FE74", x"FE69", x"FE6A", x"FE88", x"FE9F", x"FEBA", x"FED3", x"FEF5", x"FF0E", x"FF3C", x"FF6B", x"FFA3", x"FFD4", x"0010", x"0042", x"005B", x"006D", x"006C", x"0066", x"0051", x"004A", x"002B", x"0007", x"FFDA", x"FFB1", x"FF8F", x"FF7C", x"FF79", x"FF75", x"FF71", x"FF6B", x"FF6B", x"FF66", x"FF67", x"FF6F", x"FF73", x"FF80", x"FF8B", x"FF9F", x"FFA5", x"FFB0", x"FFAA", x"FFA4", x"FF98", x"FF84", x"FF7C", x"FF6A", x"FF63", x"FF5A", x"FF4C", x"FF2F", x"FF04", x"FED9", x"FEAA", x"FE83", x"FE64", x"FE55", x"FE4A", x"FE49", x"FE52", x"FE58", x"FE4D", x"FE4B", x"FE42", x"FE39", x"FE38", x"FE3E", x"FE34", x"FE26", x"FE1F", x"FE16", x"FE18", x"FE24", x"FE31", x"FE3D", x"FE3D", x"FE46", x"FE4D", x"FE58", x"FE73", x"FE95", x"FEB1", x"FEDF", x"FEF7", x"FF1C", x"FF26", x"FF3D", x"FF3B", x"FF39", x"FF2A", x"FF13", x"FEFD", x"FEE3", x"FEDA", x"FED1", x"FED4", x"FEC9", x"FEBD", x"FEB4", x"FEA1", x"FE9B", x"FE99", x"FE9A", x"FE99", x"FEA4", x"FEA8", x"FEB3", x"FEB0", x"FEB0", x"FEAA", x"FE9B", x"FE9C", x"FE93", x"FE7E", x"FE67", x"FE49", x"FE25", x"FE0E", x"FE06", x"FE00", x"FDF7", x"FDED", x"FDDC", x"FDCA", x"FDBA", x"FDB6", x"FDB3", x"FDB9", x"FDC5", x"FDDC", x"FDF8", x"FE1D", x"FE41", x"FE68", x"FE83", x"FE9B", x"FEA5", x"FEA7", x"FEA3", x"FE94", x"FE93", x"FE7E", x"FE6E", x"FE4C", x"FE2E", x"FE06", x"FDF0", x"FDE7", x"FDE2", x"FDEF", x"FE05", x"FE1D", x"FE39", x"FE49", x"FE5C", x"FE66", x"FE6E", x"FE88", x"FE92", x"FE9F", x"FE9F", x"FEA1", x"FE90", x"FE89", x"FE82", x"FE6F", x"FE5D", x"FE43", x"FE3A", x"FE32", x"FE37", x"FE4E", x"FE64", x"FE83", x"FEA2", x"FEC5", x"FEDC", x"FEE3", x"FEEF", x"FEDD", x"FECD", x"FEB9", x"FE94", x"FE74", x"FE49", x"FE34", x"FE27", x"FE19", x"FE17", x"FE05", x"FDF9", x"FDEB", x"FDF4", x"FE00", x"FE16", x"FE2C", x"FE45", x"FE4E", x"FE59", x"FE53", x"FE50", x"FE43", x"FE40", x"FE44", x"FE3B", x"FE30", x"FE12", x"FDF4", x"FDD2", x"FDB7", x"FDAA", x"FD9A", x"FD86", x"FD7B", x"FD6F", x"FD64", x"FD65", x"FD6A", x"FD6C", x"FD72", x"FD89", x"FD9B", x"FDB9", x"FDD6", x"FDF4", x"FE07", x"FE1C", x"FE26", x"FE32", x"FE32", x"FE41", x"FE51", x"FE62", x"FE7B", x"FE85", x"FE8A", x"FE7E", x"FE70", x"FE58", x"FE45", x"FE2F", x"FE1D", x"FE17", x"FE08", x"FDF9", x"FDF1", x"FDE3", x"FDE3", x"FDEA", x"FE01", x"FE0D", x"FE1C", x"FE2D", x"FE39", x"FE4B", x"FE61", x"FE7C", x"FE88", x"FE95", x"FEA3", x"FEB1", x"FEC0", x"FEDF", x"FEFB", x"FF11", x"FF2C", x"FF48", x"FF54", x"FF62", x"FF5F", x"FF58", x"FF46", x"FF3A", x"FF30", x"FF21", x"FF1B", x"FF1B", x"FF21", x"FF2C", x"FF34", x"FF37", x"FF27", x"FF12", x"FEFB", x"FEEC", x"FED8", x"FED3", x"FEC6", x"FEC0", x"FEB5", x"FEAA", x"FEA2", x"FE8B", x"FE84", x"FE7D", x"FE7F", x"FE82", x"FE85", x"FE84", x"FE6E", x"FE6D", x"FE60", x"FE67", x"FE67", x"FE75", x"FE81", x"FE8D", x"FEA1", x"FEB5", x"FEBE", x"FEC1", x"FECA", x"FED2", x"FEDC", x"FEF4", x"FF04", x"FF1D", x"FF2E", x"FF44", x"FF50", x"FF4C", x"FF48", x"FF3C", x"FF38", x"FF32", x"FF2F", x"FF28", x"FF0D", x"FEF8", x"FEE0", x"FECF", x"FEC6", x"FEC0", x"FEC3", x"FEC3", x"FEC8", x"FECD", x"FED1", x"FECE", x"FED3", x"FEE2", x"FEEE", x"FEF8", x"FF02", x"FEFE", x"FEFD", x"FEF7", x"FEFB", x"FEFA", x"FEF3", x"FEF6", x"FEF5", x"FEFD", x"FF0C", x"FF22", x"FF2B", x"FF38", x"FF4E", x"FF5E", x"FF6A", x"FF6B", x"FF63", x"FF49", x"FF2D", x"FF1C", x"FF04", x"FEE7", x"FEDE", x"FEDF", x"FEF0", x"FF13", x"FF38", x"FF53", x"FF67", x"FF7C", x"FF9E", x"FFC6", x"0002", x"0044", x"0082", x"00B9", x"00E1", x"00FF", x"0104", x"0103", x"00F8", x"00EE", x"00D9", x"00C0", x"00A0", x"0076", x"0050", x"002E", x"001A", x"FFFA", x"FFF2", x"FFE9", x"FFE8", x"FFEA", x"FFF4", x"FFF8", x"FFF7", x"FFF6", x"FFFB", x"FFFD", x"000B", x"0019", x"002A", x"0034", x"0046", x"0055", x"0058", x"005C", x"005C", x"0059", x"0053", x"0055", x"004F", x"0046", x"003B", x"0031", x"001F", x"0021", x"0016", x"001C", x"0015", x"0012", x"0006", x"FFF7", x"FFE4", x"FFD4", x"FFD1", x"FFD5", x"FFDA", x"FFE6", x"FFF2", x"FFF9", x"0005", x"0019", x"0027", x"003C", x"004B", x"0063", x"006B", x"0089", x"009E", x"00B9", x"00CB", x"00DE", x"00FE", x"010D", x"012E", x"0142", x"0143", x"013E", x"012D", x"0119", x"00FA", x"00E2", x"00D1", x"00C4", x"00CA", x"00D8", x"00E3", x"00EC", x"00E3", x"00E8", x"00DD", x"00EA", x"00F5", x"010E", x"0116", x"0126", x"0128", x"0122", x"0114", x"0109", x"0101", x"00F7", x"00F6", x"00F8", x"00E9", x"00D9", x"00C7", x"00B6", x"00A9", x"009F", x"009A", x"008B", x"0081", x"0085", x"0088", x"0091", x"00A0", x"00AE", x"00C9", x"00DA", x"0101", x"0119", x"0136", x"0150", x"016B", x"017E", x"0185", x"018B", x"0187", x"018C", x"018C", x"0199", x"018F", x"0181", x"016D", x"015A", x"014E", x"0159", x"0169", x"0181", x"0192", x"01AB", x"01B7", x"01C4", x"01D1", x"01E3", x"01FC", x"021B", x"0242", x"0255", x"0261", x"025B", x"0256", x"0243", x"023B", x"0227", x"021D", x"0205", x"0200", x"01F3", x"01FB", x"01F8", x"0203", x"0213", x"0228", x"023C", x"0255", x"025C", x"025A", x"024D", x"0241", x"0224", x"020D", x"01F4", x"01E2", x"01DA", x"01E0", x"01F1", x"01EE", x"01F0", x"01E3", x"01DF", x"01D8", x"01E8", x"01F6", x"0208", x"0218", x"0223", x"022A", x"022B", x"0233", x"0232", x"0233", x"0230", x"0220", x"020E", x"01E6", x"01CB", x"01A7", x"0192", x"0180", x"0176", x"016C", x"016D", x"016A", x"0174", x"017B", x"0185", x"019B", x"01AF", x"01C7", x"01DF", x"01FB", x"0209", x"021B", x"0229", x"0237", x"0241", x"024B", x"0257", x"0255", x"0264", x"0269", x"0275", x"026D", x"0263", x"024B", x"0229", x"0215", x"0204", x"01FD", x"01EF", x"01EB", x"01D8", x"01C8", x"01B4", x"01B1", x"01AB", x"01BC", x"01CF", x"01EB", x"01FB", x"0211", x"0217", x"0229", x"0235", x"024A", x"0261", x"026F", x"027B", x"028B", x"0298", x"02AC", x"02BD", x"02D0", x"02D5", x"02E0", x"02E7", x"02ED", x"02EE", x"02F4", x"02F3", x"02F5", x"02F1", x"02E9", x"02DD", x"02D0", x"02C9", x"02CE", x"02C9", x"02C2", x"02B5", x"0293", x"027F", x"026D", x"0267", x"0268", x"0260", x"0263", x"024A", x"023B", x"0222", x"0216", x"0207", x"020B", x"0214", x"021A", x"021E", x"021C", x"021D", x"0223", x"0231", x"0248", x"025B", x"0269", x"0271", x"0275", x"0270", x"026D", x"0264", x"0260", x"0252", x"024E", x"0246", x"024A", x"0243", x"024E", x"024D", x"024C", x"0247", x"0242", x"0234", x"0232", x"0234", x"023C", x"0231", x"0222", x"0203", x"01DC", x"01BD", x"01AD", x"01A8", x"01A5", x"01A0", x"019C", x"0183", x"0175", x"0167", x"015C", x"015C", x"0169", x"0176", x"0189", x"0191", x"01A0", x"01A1", x"019F", x"01A5", x"01A0", x"0197", x"0188", x"017A", x"0165", x"015C", x"0156", x"015B", x"0168", x"0172", x"018A", x"0191", x"01A2", x"0197", x"01A0", x"018F", x"0185", x"017E", x"016E", x"0166", x"0165", x"0177", x"0186", x"0199", x"01B1", x"01BA", x"01CC", x"01E7", x"0212", x"0242", x"026F", x"029F", x"02B0", x"02B9", x"02BC", x"02B9", x"02B0", x"02AE", x"02A1", x"028C", x"026A", x"0245", x"021A", x"01F7", x"01E1", x"01CD", x"01CC", x"01C3", x"01BF", x"01B9", x"01B3", x"01AF", x"01AD", x"01B1", x"01B5", x"01B4", x"01BB", x"01BB", x"01B9", x"01B9", x"01BD", x"01BE", x"01BF", x"01B9", x"01AE", x"0193", x"0190", x"0187", x"018C", x"018F", x"0190", x"0177", x"0163", x"0147", x"013B", x"012D", x"012A", x"0120", x"010B", x"00F2", x"00DC", x"00CA", x"00BE", x"00C1", x"00C5", x"00CA", x"00CA", x"00CF", x"00CD", x"00D5", x"00DE", x"00F0", x"00FC", x"0105", x"010A", x"0117", x"0129", x"0147", x"0175", x"0196", x"01BC", x"01D1", x"01E4", x"01EC", x"01E0", x"01E0", x"01C1", x"01A7", x"0184", x"015A", x"0132", x"010C", x"00FF", x"00F2", x"00F1", x"00FB", x"00EB", x"00E5", x"00CD", x"00D3", x"00D1", x"00E1", x"00F0", x"00F1", x"00E7", x"00D1", x"00BA", x"00A0", x"0095", x"0088", x"008B", x"007C", x"007B", x"0067", x"0060", x"0056", x"0052", x"0050", x"0047", x"003C", x"0031", x"002E", x"0027", x"002D", x"002D", x"0031", x"002D", x"002E", x"0034", x"0038", x"0049", x"0061", x"0072", x"0087", x"0093", x"0095", x"0095", x"0095", x"00A1", x"00A4", x"00B0", x"00A8", x"0093", x"0074", x"0056", x"0049", x"0044", x"0053", x"0062", x"006E", x"0071", x"0072", x"0071", x"0070", x"0077", x"008B", x"0092", x"009B", x"0094", x"008C", x"007A", x"006F", x"0069", x"0062", x"0058", x"004A", x"0039", x"0025", x"001C", x"001B", x"002F", x"0041", x"005F", x"0075", x"0088", x"008C", x"008C", x"0084", x"0069", x"0057", x"0035", x"0018", x"FFF5", x"FFE4", x"FFD6", x"FFD7", x"FFDF", x"FFED", x"FFE5", x"FFE7", x"FFE3", x"FFEF", x"FFFE", x"001F", x"0036", x"0046", x"0042", x"003A", x"0026", x"0018", x"0011", x"FFFE", x"FFEC", x"FFC8", x"FF9D", x"FF6E", x"FF43", x"FF23", x"FF05", x"FEEF", x"FED5", x"FEB5", x"FE9B", x"FE7E", x"FE72", x"FE71", x"FE81", x"FE8C", x"FEA2", x"FEB6", x"FECB", x"FEE7", x"FF0B", x"FF35", x"FF5A", x"FF7B", x"FF8F", x"FF92", x"FF86", x"FF86", x"FF75", x"FF6F", x"FF66", x"FF51", x"FF33", x"FF0C", x"FEEB", x"FECD", x"FEC2", x"FEB5", x"FEB3", x"FE9D", x"FE8E", x"FE76", x"FE67", x"FE67", x"FE6F", x"FE7C", x"FE8B", x"FE94", x"FE9C", x"FEA3", x"FEB2", x"FEC6", x"FEDE", x"FEEE", x"FEEE", x"FEEC", x"FEE1", x"FEDF", x"FEE4", x"FEF9", x"FF09", x"FF1B", x"FF24", x"FF2A", x"FF2B", x"FF34", x"FF41", x"FF44", x"FF50", x"FF42", x"FF37", x"FF18", x"FF00", x"FEF0", x"FEE4", x"FEEA", x"FEF1", x"FEF7", x"FEF3", x"FEED", x"FEE8", x"FEE2", x"FEF6", x"FEF6", x"FF00", x"FEF3", x"FED6", x"FEB2", x"FE8D", x"FE6E", x"FE5F", x"FE57", x"FE5B", x"FE60", x"FE65", x"FE6D", x"FE75", x"FE80", x"FE8D", x"FE91", x"FE95", x"FE88", x"FE82", x"FE6B", x"FE66", x"FE5D", x"FE5C", x"FE56", x"FE4F", x"FE49", x"FE41", x"FE4A", x"FE4C", x"FE5F", x"FE61", x"FE66", x"FE56", x"FE4A", x"FE39", x"FE31", x"FE35", x"FE30", x"FE2F", x"FE20", x"FE04", x"FDEB", x"FDCF", x"FDCA", x"FDC8", x"FDD6", x"FDDF", x"FDDE", x"FDD3", x"FDC4", x"FDB7", x"FDBB", x"FDC7", x"FDDE", x"FDF6", x"FE05", x"FE0E", x"FE0F", x"FE13", x"FE15", x"FE19", x"FE1B", x"FE11", x"FE01", x"FDE9", x"FDD9", x"FDD2", x"FDD9", x"FDEA", x"FDF8", x"FE03", x"FE05", x"FE01", x"FE00", x"FDFB", x"FDFC", x"FDF6", x"FDEC", x"FDDC", x"FDD4", x"FDD0", x"FDE3", x"FDFB", x"FE24", x"FE47", x"FE66", x"FE80", x"FE9B", x"FEBD", x"FEE9", x"FF19", x"FF42", x"FF56", x"FF57", x"FF46", x"FF2E", x"FF13", x"FF01", x"FEEB", x"FED0", x"FEB2", x"FE8A", x"FE5E", x"FE3A", x"FE20", x"FE10", x"FE0E", x"FE05", x"FDFD", x"FDF0", x"FDDE", x"FDDD", x"FDD8", x"FDEC", x"FDF5", x"FDFC", x"FE02", x"FE00", x"FE01", x"FE11", x"FE23", x"FE3A", x"FE4B", x"FE4A", x"FE41", x"FE2B", x"FE1E", x"FE17", x"FE16", x"FE19", x"FE17", x"FE0E", x"FDFB", x"FDEC", x"FDE1", x"FDE3", x"FDEA", x"FDF3", x"FDF5", x"FDEC", x"FDDF", x"FDD1", x"FDC9", x"FDCC", x"FDD1", x"FDDD", x"FDE9", x"FDEC", x"FDFB", x"FDFF", x"FE11", x"FE1C", x"FE2A", x"FE2D", x"FE2C", x"FE27", x"FE29", x"FE2B", x"FE4A", x"FE67", x"FE92", x"FEAD", x"FEC3", x"FECA", x"FEC7", x"FEC9", x"FEC9", x"FECC", x"FEBD", x"FEB1", x"FE89", x"FE6D", x"FE4A", x"FE43", x"FE3C", x"FE4C", x"FE53", x"FE5C", x"FE5F", x"FE6A", x"FE7B", x"FE97", x"FEBC", x"FED5", x"FEE3", x"FED9", x"FEB8", x"FE99", x"FE6B", x"FE56", x"FE41", x"FE42", x"FE45", x"FE49", x"FE54", x"FE56", x"FE5E", x"FE63", x"FE67", x"FE69", x"FE61", x"FE54", x"FE4A", x"FE3E", x"FE3E", x"FE48", x"FE4C", x"FE56", x"FE5A", x"FE64", x"FE71", x"FE91", x"FEB9", x"FED5", x"FEF0", x"FEF1", x"FEE6", x"FED4", x"FECD", x"FECA", x"FECE", x"FECF", x"FEC9", x"FEB7", x"FEA2", x"FE9C", x"FEAB", x"FECC", x"FEFC", x"FF24", x"FF3D", x"FF47", x"FF3F", x"FF41", x"FF3C", x"FF4C", x"FF4F", x"FF5E", x"FF5B", x"FF55", x"FF4B", x"FF45", x"FF3A", x"FF37", x"FF2C", x"FF16", x"FEEE", x"FECD", x"FEA0", x"FE8C", x"FE8E", x"FEA4", x"FEC2", x"FEDF", x"FEFE", x"FF0A", x"FF1E", x"FF2E", x"FF3E", x"FF42", x"FF42", x"FF29", x"FF13", x"FEF6", x"FEEE", x"FEEB", x"FEF3", x"FEFE", x"FEFB", x"FEF2", x"FEEB", x"FEEB", x"FEF6", x"FF17", x"FF2F", x"FF40", x"FF3E", x"FF31", x"FF11", x"FEFE", x"FEE8", x"FEDE", x"FED9", x"FEDB", x"FED6", x"FED4", x"FECA", x"FECB", x"FEBC", x"FEBE", x"FEB3", x"FEA8", x"FE8F", x"FE7B", x"FE63", x"FE60", x"FE69", x"FE81", x"FE9B", x"FEC0", x"FED9", x"FEF6", x"FF1A", x"FF3E", x"FF69", x"FF93", x"FFB7", x"FFBF", x"FFC1", x"FFB3", x"FFA8", x"FF9E", x"FF97", x"FF90", x"FF79", x"FF68", x"FF54", x"FF44", x"FF47", x"FF52", x"FF5A", x"FF65", x"FF61", x"FF5E", x"FF4B", x"FF49", x"FF40", x"FF4B", x"FF53", x"FF5F", x"FF69", x"FF70", x"FF7A", x"FF85", x"FF91", x"FFAC", x"FFAF", x"FFBB", x"FFBA", x"FFB8", x"FFB6", x"FFC6", x"FFDB", x"FFF6", x"0012", x"0028", x"002B", x"0032", x"0031", x"003F", x"0043", x"004F", x"0047", x"002D", x"0011", x"FFF9", x"FFED", x"FFF0", x"0004", x"000B", x"000E", x"0004", x"FFFB", x"FFFC", x"0007", x"0025", x"0036", x"0046", x"0039", x"0021", x"FFFE", x"FFE5", x"FFD5", x"FFE1", x"FFF3", x"001B", x"0038", x"0064", x"0085", x"00AB", x"00CA", x"00E8", x"00F1", x"00EB", x"00D7", x"00B8", x"0095", x"007F", x"0069", x"0061", x"0053", x"0049", x"003A", x"0033", x"0036", x"0045", x"0054", x"0068", x"0065", x"0065", x"0055", x"0053", x"0052", x"0058", x"0057", x"004E", x"0031", x"001B", x"0004", x"0002", x"000D", x"0027", x"0030", x"003C", x"0024", x"0013", x"FFEC", x"FFE5", x"FFD2", x"FFE4", x"FFED", x"FFFE", x"0008", x"000F", x"0015", x"001C", x"002B", x"0035", x"0038", x"0035", x"0027", x"0016", x"000E", x"000F", x"0019", x"002B", x"0041", x"0054", x"0060", x"006D", x"007C", x"0083", x"0096", x"009C", x"00A2", x"009B", x"009D", x"00A0", x"00AC", x"00CA", x"00DD", x"00F5", x"0103", x"0118", x"012B", x"014E", x"017A", x"01A7", x"01C3", x"01DF", x"01D8", x"01CB", x"01B5", x"01A1", x"018B", x"0181", x"0175", x"016D", x"015C", x"014D", x"0140", x"0133", x"012E", x"0130", x"0121", x"0112", x"00FA", x"00DF", x"00D3", x"00CF", x"00DF", x"00F3", x"0114", x"0125", x"013B", x"0151", x"015E", x"017D", x"018F", x"01A0", x"0198", x"018D", x"0171", x"015F", x"014B", x"014A", x"0135", x"012A", x"0117", x"0109", x"010A", x"0117", x"0137", x"0153", x"0166", x"0171", x"015E", x"0148", x"0128", x"0116", x"010F", x"0115", x"0123", x"0130", x"0139", x"0144", x"0152", x"016B", x"017B", x"0187", x"0189", x"0182", x"0173", x"017A", x"0187", x"01A9", x"01D0", x"01FD", x"021E", x"022F", x"0235", x"023A", x"022F", x"0231", x"0226", x"020F", x"01E4", x"01BF", x"0193", x"017B", x"0179", x"017D", x"018A", x"0190", x"019A", x"01AA", x"01C1", x"01EF", x"0225", x"0256", x"027A", x"0281", x"026F", x"024B", x"0220", x"01FE", x"01E5", x"01D9", x"01D4", x"01CF", x"01CB", x"01CA", x"01C6", x"01CD", x"01CC", x"01C8", x"01BD", x"01A0", x"0189", x"016A", x"015C", x"0155", x"015D", x"0168", x"017D", x"0186", x"019D", x"01AD", x"01C7", x"01DA", x"01F0", x"01FC", x"0201", x"0206", x"0208", x"020E", x"0211", x"020F", x"0205", x"01EC", x"01DC", x"01D1", x"01D7", x"01F0", x"0212", x"0235", x"024B", x"0252", x"024D", x"022E", x"0227", x"020D", x"0213", x"0216", x"0223", x"022A", x"022D", x"0234", x"023F", x"024D", x"0258", x"0256", x"0248", x"0223", x"0209", x"01E8", x"01E0", x"01E5", x"01FE", x"021A", x"023C", x"0250", x"0268", x"026A", x"0274", x"0273", x"027A", x"026C", x"0263", x"0251", x"023D", x"0239", x"0237", x"0236", x"0229", x"021D", x"0209", x"0205", x"0206", x"0225", x"023B", x"0256", x"025E", x"025C", x"023D", x"022D", x"020D", x"0202", x"01FB", x"0200", x"01F6", x"01F1", x"01DC", x"01CD", x"01BE", x"01B0", x"01AA", x"018E", x"016E", x"0142", x"0115", x"00FE", x"00F8", x"010C", x"012B", x"0159", x"017A", x"01A5", x"01C5", x"01EA", x"0215", x"023A", x"0265", x"026F", x"0279", x"026A", x"0253", x"023F", x"0220", x"01F6", x"01C4", x"0193", x"0163", x"014D", x"0148", x"015B", x"0172", x"0188", x"019E", x"019A", x"0191", x"0186", x"017D", x"017D", x"0185", x"0191", x"0197", x"0199", x"0198", x"01A4", x"01AC", x"01BB", x"01C1", x"01BB", x"01A7", x"018E", x"0180", x"0175", x"017A", x"018D", x"01A6", x"01BC", x"01CD", x"01DC", x"01DB", x"01D7", x"01D4", x"01CE", x"01C0", x"01AB", x"0199", x"0181", x"017C", x"0177", x"0186", x"017E", x"0182", x"017D", x"017F", x"0188", x"01A7", x"01CB", x"01EE", x"0204", x"020C", x"01F7", x"01DA", x"01B1", x"0190", x"0174", x"016E", x"016C", x"0173", x"0184", x"018C", x"01A5", x"01AD", x"01C2", x"01C2", x"01B8", x"01A0", x"0175", x"014E", x"0131", x"011A", x"011E", x"0121", x"0135", x"0134", x"013D", x"013B", x"0136", x"0136", x"0132", x"012C", x"0123", x"0118", x"0113", x"0101", x"00FA", x"00E7", x"00CA", x"00AD", x"0094", x"0082", x"0081", x"0095", x"00B4", x"00CC", x"00DC", x"00DB", x"00BE", x"00A0", x"007F", x"0064", x"005D", x"005D", x"0060", x"0068", x"0067", x"0075", x"007C", x"0097", x"00A5", x"00B6", x"00A9", x"0096", x"006E", x"0050", x"0032", x"002B", x"002C", x"0039", x"0044", x"0055", x"005B", x"0064", x"006C", x"007E", x"008F", x"0099", x"00AD", x"00B0", x"00B9", x"00CD", x"00E9", x"00FD", x"010C", x"0112", x"010C", x"0108", x"0118", x"0129", x"013D", x"0148", x"014D", x"0136", x"011F", x"0104", x"00E4", x"00CE", x"00BC", x"00B5", x"00A3", x"0098", x"008C", x"0079", x"0077", x"0070", x"006D", x"0054", x"003D", x"0005", x"FFDC", x"FFAD", x"FF9A", x"FF92", x"FFA3", x"FFB8", x"FFCF", x"FFE1", x"FFF0", x"FFF8", x"0003", x"0011", x"0015", x"001C", x"0016", x"0010", x"FFFC", x"FFED", x"FFD5", x"FFB4", x"FF95", x"FF78", x"FF64", x"FF63", x"FF7F", x"FF9C", x"FFC6", x"FFE5", x"FFFB", x"FFFA", x"FFF0", x"FFDB", x"FFC7", x"FFB4", x"FFAF", x"FFAD", x"FFAF", x"FFB4", x"FFBB", x"FFC1", x"FFCD", x"FFD1", x"FFD1", x"FFC2", x"FFA9", x"FF90", x"FF7A", x"FF6F", x"FF69", x"FF7D", x"FF8E", x"FFAA", x"FFBB", x"FFCD", x"FFC7", x"FFBB", x"FFB5", x"FFA3", x"FF90", x"FF81", x"FF63", x"FF46", x"FF2E", x"FF26", x"FF23", x"FF1A", x"FF22", x"FF14", x"FF18", x"FF2C", x"FF4D", x"FF74", x"FF9C", x"FFB5", x"FFBA", x"FFB0", x"FF98", x"FF7A", x"FF57", x"FF36", x"FF2A", x"FF0F", x"FF11", x"FF05", x"FF06", x"FF03", x"FF0D", x"FF0E", x"FF14", x"FF09", x"FEEE", x"FEC5", x"FE9F", x"FE7E", x"FE74", x"FE79", x"FE96", x"FEAE", x"FEC9", x"FED6", x"FEE2", x"FEE1", x"FEF5", x"FEF9", x"FF07", x"FF10", x"FF16", x"FF18", x"FF1E", x"FF21", x"FF1C", x"FF0F", x"FEFD", x"FEE8", x"FEE1", x"FEEE", x"FF10", x"FF3D", x"FF71", x"FF96", x"FFA3", x"FFA3", x"FF8E", x"FF75", x"FF54", x"FF42", x"FF27", x"FF19", x"FF09", x"FF01", x"FEF8", x"FF00", x"FF07", x"FF0B", x"FF09", x"FEF3", x"FED3", x"FEA6", x"FE88", x"FE63", x"FE60", x"FE64", x"FE7B", x"FE91", x"FEB1", x"FEB8", x"FEC2", x"FEC0", x"FEC8", x"FEC1", x"FEC7", x"FEBF", x"FEB5", x"FEA2", x"FEA3", x"FE96", x"FE92", x"FE83", x"FE76", x"FE58", x"FE51", x"FE5F", x"FE69", x"FE87", x"FE94", x"FE99", x"FE87", x"FE7E", x"FE69", x"FE5A", x"FE44", x"FE40", x"FE31", x"FE2C", x"FE2E", x"FE2E", x"FE30", x"FE39", x"FE3F", x"FE3A", x"FE31", x"FE16", x"FDF5", x"FDCA", x"FDAA", x"FD8D", x"FD90", x"FD9B", x"FDBC", x"FDD3", x"FDF7", x"FE09", x"FE1F", x"FE35", x"FE50", x"FE69", x"FE84", x"FE93", x"FE98", x"FE90", x"FE89", x"FE70", x"FE4A", x"FE30", x"FDFC", x"FDDF", x"FDCC", x"FDD6", x"FDE5", x"FE0E", x"FE29", x"FE3F", x"FE3E", x"FE3F", x"FE28", x"FE13", x"FE02", x"FDF4", x"FDE9", x"FDE9", x"FDEC", x"FDF4", x"FE00", x"FE13", x"FE22", x"FE30", x"FE33", x"FE2C", x"FE18", x"FE06", x"FDF8", x"FDED", x"FE02", x"FE15", x"FE37", x"FE51", x"FE69", x"FE66", x"FE67", x"FE62", x"FE58", x"FE55", x"FE50", x"FE3B", x"FE2A", x"FE19", x"FE16", x"FE0B", x"FE0C", x"FE05", x"FDF4", x"FDE9", x"FDF2", x"FE0F", x"FE34", x"FE68", x"FE91", x"FEA2", x"FEA3", x"FEA2", x"FE86", x"FE7A", x"FE6E", x"FE6C", x"FE6F", x"FE87", x"FE9A", x"FEB6", x"FED0", x"FEE5", x"FEF5", x"FEF3", x"FEE5", x"FEBB", x"FE88", x"FE52", x"FE1A", x"FE00", x"FDF0", x"FDFD", x"FE02", x"FE1C", x"FE1D", x"FE19", x"FE1B", x"FE1A", x"FE1F", x"FE2B", x"FE37", x"FE37", x"FE31", x"FE31", x"FE22", x"FE14", x"FDFB", x"FDDD", x"FDB4", x"FD9A", x"FDA1", x"FDA8", x"FDD0", x"FDF3", x"FE0C", x"FE0F", x"FE10", x"FDFA", x"FDE8", x"FDCB", x"FDBE", x"FD9F", x"FD97", x"FD97", x"FD98", x"FDAE", x"FDC5", x"FDE4", x"FE02", x"FE14", x"FE20", x"FE10", x"FE00", x"FDE5", x"FDCE", x"FDC3", x"FDCA", x"FDD2", x"FDF4", x"FE09", x"FE23", x"FE30", x"FE3E", x"FE46", x"FE51", x"FE5E", x"FE6C", x"FE6D", x"FE72", x"FE80", x"FE82", x"FE95", x"FEA2", x"FEA2", x"FE96", x"FE96", x"FE99", x"FEA9", x"FEC6", x"FEE5", x"FEF6", x"FEFC", x"FF01", x"FEF3", x"FEE5", x"FEDD", x"FED1", x"FEC9", x"FEC5", x"FEC4", x"FEC5", x"FECA", x"FECC", x"FECF", x"FEC3", x"FEB5", x"FE8C", x"FE64", x"FE36", x"FE08", x"FDF2", x"FDEB", x"FDFB", x"FE15", x"FE3E", x"FE59", x"FE6C", x"FE74", x"FE88", x"FE91", x"FEA7", x"FEC4", x"FECB", x"FEC5", x"FEBC", x"FEAF", x"FE92", x"FE88", x"FE71", x"FE5A", x"FE41", x"FE3A", x"FE43", x"FE5A", x"FE8A", x"FEB5", x"FED0", x"FEE3", x"FEE2", x"FED7", x"FEC3", x"FEB8", x"FEB4", x"FEAC", x"FEBF", x"FEC5", x"FED7", x"FEE5", x"FEF6", x"FF06", x"FF11", x"FF1C", x"FF0A", x"FF03", x"FEE5", x"FED2", x"FEC6", x"FECD", x"FED6", x"FEEC", x"FEFE", x"FF0D", x"FF09", x"FF09", x"FF02", x"FEF5", x"FEF6", x"FEF6", x"FEEE", x"FEEE", x"FEF6", x"FEF8", x"FF0D", x"FF1B", x"FF2C", x"FF28", x"FF2C", x"FF3A", x"FF48", x"FF74", x"FFA0", x"FFC8", x"FFD7", x"FFDF", x"FFCA", x"FFAE", x"FF91", x"FF73", x"FF5A", x"FF47", x"FF3F", x"FF3E", x"FF45", x"FF5D", x"FF68", x"FF7B", x"FF7E", x"FF70", x"FF52", x"FF32", x"FF0B", x"FEEB", x"FEE5", x"FEE9", x"FF00", x"FF23", x"FF4C", x"FF5C", x"FF70", x"FF70", x"FF7C", x"FF7F", x"FF9D", x"FFBB", x"FFC9", x"FFE2", x"FFF0", x"FFFF", x"0001", x"0014", x"0003", x"FFF3", x"FFE4", x"FFE2", x"FFE7", x"000A", x"0025", x"0046", x"0049", x"004C", x"0034", x"0015", x"FFF5", x"FFD1", x"FFB9", x"FFA7", x"FFAA", x"FFB0", x"FFCE", x"FFEF", x"0019", x"0042", x"0062", x"0071", x"0069", x"005B", x"0037", x"001E", x"000B", x"0006", x"0013", x"002F", x"004D", x"005D", x"0073", x"0073", x"007E", x"0087", x"009E", x"00AB", x"00B4", x"00BE", x"00BC", x"00BC", x"00C3", x"00C9", x"00C0", x"00B4", x"00A4", x"008F", x"0089", x"0097", x"00A7", x"00B8", x"00C4", x"00C2", x"00B1", x"009C", x"0089", x"0076", x"0066", x"0064", x"0058", x"0060", x"0067", x"0073", x"0081", x"0085", x"0084", x"006A", x"004F", x"002C", x"000C", x"FFF5", x"FFF4", x"FFF9", x"0012", x"0038", x"0057", x"0070", x"0086", x"009E", x"00A9", x"00CE", x"00E5", x"00F8", x"00FC", x"00F6", x"00F0", x"00DD", x"00D8", x"00C8", x"00AF", x"0098", x"0086", x"0087", x"0091", x"00C1", x"00E5", x"010C", x"0124", x"0125", x"011C", x"0103", x"00E7", x"00CF", x"00B7", x"00AE", x"00A3", x"00A8", x"00AE", x"00C0", x"00D1", x"00E5", x"00ED", x"00EB", x"00EA", x"00DB", x"00D7", x"00DB", x"00E6", x"0106", x"0122", x"014E", x"0163", x"0177", x"0181", x"017A", x"0175", x"0173", x"016B", x"0163", x"015B", x"0152", x"014F", x"014D", x"0158", x"0158", x"0157", x"015C", x"0165", x"0178", x"01A3", x"01D2", x"01F9", x"0219", x"0220", x"0211", x"01F2", x"01D0", x"01AF", x"0192", x"0185", x"0184", x"0185", x"0199", x"01AC", x"01BC", x"01D0", x"01D7", x"01D3", x"01C5", x"01B2", x"0197", x"0182", x"017B", x"017B", x"018B", x"01A6", x"01C2", x"01CF", x"01CE", x"01C7", x"01B0", x"01A5", x"01A0", x"01A1", x"0194", x"018F", x"017F", x"0173", x"0169", x"0164", x"0159", x"0142", x"013D", x"0130", x"0139", x"0152", x"0177", x"0195", x"01B6", x"01BE", x"01BF", x"01A3", x"018B", x"0168", x"014B", x"0139", x"0129", x"012F", x"013B", x"0159", x"017D", x"01A8", x"01C2", x"01D4", x"01D1", x"01C6", x"01AA", x"0199", x"0189", x"018E", x"0196", x"01BE", x"01D1", x"01EA", x"01F3", x"01FB", x"01FE", x"020D", x"0221", x"0231", x"023E", x"024C", x"0252", x"025D", x"0264", x"0266", x"025A", x"0246", x"0231", x"0220", x"021A", x"022B", x"0239", x"0251", x"0262", x"0261", x"025D", x"024A", x"0240", x"022A", x"0229", x"021F", x"0222", x"0221", x"0230", x"0233", x"0239", x"022F", x"0219", x"01EF", x"01BE", x"0186", x"0153", x"012A", x"011C", x"0114", x"0126", x"013E", x"0159", x"0168", x"0181", x"0195", x"01AE", x"01CC", x"01E9", x"01F5", x"01FB", x"01FF", x"01FA", x"01F8", x"01F9", x"01EE", x"01E1", x"01C5", x"01B9", x"01A4", x"01B2", x"01C2", x"01E6", x"0203", x"0224", x"0232", x"0236", x"0230", x"0224", x"020F", x"0204", x"01F1", x"01E9", x"01E2", x"01E2", x"01E4", x"01E1", x"01E5", x"01D1", x"01C3", x"01A4", x"018B", x"015E", x"0152", x"013F", x"0148", x"015E", x"0183", x"0198", x"01AE", x"01B2", x"01B5", x"01B0", x"01B4", x"01B6", x"01AE", x"01AD", x"01A8", x"01A4", x"01A4", x"01A7", x"0198", x"018B", x"0177", x"0170", x"016F", x"0186", x"01A5", x"01CA", x"01E9", x"0208", x"0206", x"0205", x"01F4", x"01DD", x"01C8", x"01B8", x"01AB", x"01A1", x"01A3", x"01A2", x"01A7", x"01A5", x"01A5", x"018C", x"0176", x"0155", x"012D", x"010D", x"00F4", x"00EC", x"00F2", x"0109", x"0125", x"012F", x"013F", x"0143", x"0144", x"014E", x"0162", x"016D", x"017D", x"0188", x"0198", x"019F", x"01B8", x"01C9", x"01C4", x"01C8", x"01B4", x"01B1", x"01AC", x"01C1", x"01CF", x"01DE", x"01E0", x"01D3", x"01B1", x"0188", x"015C", x"0128", x"0108", x"00EA", x"00D5", x"00D4", x"00E3", x"00FC", x"012A", x"0152", x"0179", x"0189", x"018C", x"017D", x"0152", x"0136", x"0110", x"0101", x"00FD", x"010E", x"0113", x"010F", x"010B", x"00FF", x"00F8", x"0101", x"010F", x"011B", x"011E", x"012D", x"0131", x"013D", x"0149", x"014D", x"0141", x"0131", x"011A", x"0108", x"00FC", x"00FF", x"00FF", x"0107", x"0104", x"00FB", x"00E1", x"00CF", x"00AA", x"0094", x"007F", x"006D", x"005F", x"0062", x"006C", x"0071", x"008B", x"008D", x"008C", x"0078", x"0067", x"0040", x"0019", x"FFFC", x"FFE0", x"FFD4", x"FFDF", x"FFF0", x"0002", x"000D", x"0013", x"001A", x"001B", x"0039", x"004A", x"005F", x"006B", x"0078", x"0074", x"0081", x"0089", x"0084", x"0077", x"0066", x"0042", x"0034", x"002D", x"003C", x"0048", x"0063", x"0069", x"0067", x"0057", x"0045", x"0027", x"0003", x"FFEF", x"FFCA", x"FFC0", x"FFB9", x"FFC9", x"FFD3", x"FFF0", x"FFFF", x"0008", x"0002", x"0003", x"FFE5", x"FFD7", x"FFC5", x"FFC2", x"FFCA", x"FFE7", x"000A", x"001E", x"002E", x"002D", x"0027", x"001F", x"0024", x"001C", x"0016", x"0004", x"FFF9", x"FFE1", x"FFE6", x"FFE0", x"FFE1", x"FFDE", x"FFDC", x"FFD9", x"FFE3", x"FFFD", x"001A", x"0046", x"0060", x"007A", x"0070", x"006C", x"0058", x"0042", x"003D", x"0036", x"0028", x"002A", x"001C", x"001E", x"0022", x"0028", x"002A", x"0017", x"000C", x"FFE8", x"FFCA", x"FFAB", x"FF9B", x"FF85", x"FF8C", x"FF9B", x"FFA6", x"FFAB", x"FFA5", x"FF91", x"FF71", x"FF69", x"FF59", x"FF48", x"FF37", x"FF23", x"FF02", x"FEF1", x"FEE6", x"FEE6", x"FED5", x"FED7", x"FEC4", x"FEB9", x"FEBE", x"FECF", x"FEE8", x"FEFC", x"FF18", x"FF14", x"FF0D", x"FEF6", x"FEDB", x"FEB7", x"FE9F", x"FE85", x"FE71", x"FE65", x"FE6C", x"FE76", x"FE8E", x"FEB3", x"FEC5", x"FEDC", x"FEE4", x"FEE1", x"FECF", x"FEC8", x"FEBF", x"FEBE", x"FEDB", x"FEF1", x"FF11", x"FF1B", x"FF27", x"FF1D", x"FF19", x"FF23", x"FF2E", x"FF35", x"FF3E", x"FF3B", x"FF31", x"FF29", x"FF21", x"FF15", x"FF0C", x"FEFD", x"FEF5", x"FEEB", x"FEF3", x"FF00", x"FF15", x"FF2B", x"FF3E", x"FF3C", x"FF3E", x"FF2A", x"FF19", x"FF0E", x"FF01", x"FEF6", x"FEE8", x"FEE8", x"FEE2", x"FEE2", x"FEED", x"FEE6", x"FED6", x"FEBA", x"FE98", x"FE67", x"FE40", x"FE1F", x"FE07", x"FDFA", x"FE0E", x"FE22", x"FE3A", x"FE51", x"FE59", x"FE61", x"FE6A", x"FE8E", x"FEA4", x"FEC3", x"FED4", x"FEDF", x"FED4", x"FED5", x"FED3", x"FEC7", x"FEC3", x"FEA9", x"FE95", x"FE75", x"FE78", x"FE77", x"FE8D", x"FEA4", x"FEBC", x"FEC0", x"FEC3", x"FEBF", x"FEAE", x"FEAC", x"FEA7", x"FEA2", x"FE9E", x"FE9D", x"FE9C", x"FE9D", x"FEA7", x"FEAA", x"FEA5", x"FE98", x"FE75", x"FE51", x"FE1F", x"FE03", x"FDE4", x"FDEE", x"FDF1", x"FE11", x"FE1C", x"FE2E", x"FE2E", x"FE2D", x"FE2F", x"FE41", x"FE4C", x"FE61", x"FE6B", x"FE6B", x"FE69", x"FE68", x"FE6A", x"FE68", x"FE6B", x"FE63", x"FE5A", x"FE50", x"FE52", x"FE5A", x"FE6E", x"FE87", x"FE9A", x"FEA7", x"FEA9", x"FEA3", x"FE97", x"FE93", x"FE89", x"FE86", x"FE7E", x"FE7D", x"FE7C", x"FE7D", x"FE87", x"FE83", x"FE7C", x"FE6E", x"FE47", x"FE27", x"FDFD", x"FDE4", x"FDCC", x"FDCF", x"FDDD", x"FDE8", x"FDFA", x"FE01", x"FE03", x"FDFE", x"FE12", x"FE21", x"FE3C", x"FE4F", x"FE65", x"FE68", x"FE75", x"FE7D", x"FE88", x"FE82", x"FE7F", x"FE7A", x"FE67", x"FE6B", x"FE6F", x"FE71", x"FE7E", x"FE82", x"FE7D", x"FE71", x"FE57", x"FE3E", x"FE1E", x"FE08", x"FDFE", x"FDF6", x"FE00", x"FE09", x"FE25", x"FE3A", x"FE60", x"FE7E", x"FE91", x"FE9A", x"FE8F", x"FE76", x"FE5F", x"FE3F", x"FE39", x"FE39", x"FE48", x"FE59", x"FE61", x"FE6C", x"FE62", x"FE6D", x"FE7F", x"FEA4", x"FEBA", x"FEDC", x"FEE2", x"FEE4", x"FEE4", x"FEED", x"FEEE", x"FEF7", x"FEF3", x"FEE7", x"FED4", x"FEC3", x"FEB7", x"FEAD", x"FEA9", x"FEAA", x"FEA5", x"FE9F", x"FE94", x"FE85", x"FE77", x"FE74", x"FE71", x"FE75", x"FE7E", x"FE84", x"FE8F", x"FE98", x"FEA2", x"FE99", x"FE9C", x"FE86", x"FE6D", x"FE4A", x"FE2A", x"FE0C", x"FDFF", x"FE06", x"FE19", x"FE20", x"FE29", x"FE23", x"FE14", x"FE0F", x"FE2A", x"FE3B", x"FE67", x"FE81", x"FE9C", x"FEA4", x"FEB8", x"FECA", x"FECE", x"FED5", x"FECE", x"FEC1", x"FEAF", x"FEAC", x"FEA4", x"FEA9", x"FEB4", x"FEB3", x"FEB3", x"FE99", x"FE87", x"FE59", x"FE3C", x"FE18", x"FE05", x"FDF1", x"FDEF", x"FDEC", x"FDF1", x"FDFD", x"FE0F", x"FE19", x"FE26", x"FE25", x"FE21", x"FE18", x"FE18", x"FE1E", x"FE33", x"FE4F", x"FE71", x"FE88", x"FE9A", x"FE9C", x"FE96", x"FEA2", x"FEAC", x"FEC2", x"FED2", x"FED8", x"FED3", x"FEC6", x"FED0", x"FECC", x"FEE1", x"FEE5", x"FEF7", x"FEF4", x"FEFE", x"FF10", x"FF1C", x"FF31", x"FF48", x"FF52", x"FF58", x"FF5E", x"FF5A", x"FF4B", x"FF43", x"FF3C", x"FF35", x"FF38", x"FF42", x"FF44", x"FF46", x"FF51", x"FF4D", x"FF51", x"FF4D", x"FF41", x"FF29", x"FF15", x"FEFB", x"FEF2", x"FEEF", x"FF03", x"FF0A", x"FF09", x"FEFC", x"FEDD", x"FEB6", x"FEAD", x"FEA5", x"FEA5", x"FEAD", x"FEA5", x"FE99", x"FE91", x"FE9B", x"FE9E", x"FEA9", x"FEAF", x"FEB3", x"FEA5", x"FEB0", x"FEB5", x"FEBE", x"FECC", x"FEE3", x"FEE6", x"FEEB", x"FEEC", x"FEDA", x"FECA", x"FEB7", x"FEB5", x"FEAC", x"FEC1", x"FECE", x"FEE6", x"FEFA", x"FF16", x"FF27", x"FF3E", x"FF4D", x"FF57", x"FF4E", x"FF4C", x"FF41", x"FF3B", x"FF53", x"FF68", x"FF89", x"FF9E", x"FFA9", x"FF9C", x"FFA1", x"FFB0", x"FFC9", x"FFE2", x"0004", x"FFFE", x"FFF4", x"FFE5", x"FFDF", x"FFD7", x"FFD9", x"FFDF", x"FFCB", x"FFC5", x"FFC2", x"FFC7", x"FFC9", x"FFE2", x"FFEB", x"FFEC", x"FFF1", x"FFEC", x"FFE6", x"FFD4", x"FFD0", x"FFC2", x"FFBC", x"FFC9", x"FFCD", x"FFCD", x"FFCF", x"FFC4", x"FFB1", x"FF9E", x"FF8C", x"FF65", x"FF50", x"FF2E", x"FF1B", x"FF0F", x"FF24", x"FF33", x"FF4C", x"FF60", x"FF6A", x"FF72", x"FF88", x"FFB2", x"FFDB", x"0010", x"003D", x"0051", x"005A", x"0068", x"0073", x"0077", x"0086", x"007C", x"006F", x"005F", x"005F", x"005A", x"0066", x"0073", x"007C", x"007C", x"0085", x"0079", x"0072", x"0067", x"0061", x"0054", x"0054", x"004F", x"0047", x"003B", x"0036", x"0025", x"001C", x"0014", x"0005", x"FFF0", x"FFDF", x"FFCE", x"FFC5", x"FFD2", x"FFEC", x"0008", x"0027", x"003B", x"003C", x"0038", x"003A", x"0044", x"0053", x"0067", x"0070", x"005C", x"0054", x"0048", x"0046", x"004A", x"0059", x"0053", x"004B", x"004C", x"0050", x"005C", x"0079", x"009B", x"00B6", x"00D0", x"00E9", x"00F8", x"00F1", x"00FC", x"00F2", x"00F2", x"0105", x"010F", x"011C", x"011A", x"0119", x"0107", x"00F7", x"00ED", x"00D9", x"00C3", x"00AD", x"0097", x"0086", x"008C", x"0092", x"00A2", x"00A9", x"00A7", x"0093", x"0082", x"0086", x"008F", x"00B6", x"00DF", x"00FA", x"010F", x"0117", x"012A", x"012C", x"013E", x"014C", x"0140", x"0140", x"013A", x"013B", x"0137", x"0145", x"0146", x"013D", x"013A", x"0129", x"0112", x"00FE", x"00F1", x"00E2", x"00E2", x"00EC", x"00FF", x"0106", x"011E", x"0128", x"0134", x"0147", x"0152", x"0154", x"014B", x"0146", x"012A", x"0123", x"011C", x"0124", x"0124", x"0132", x"012B", x"0127", x"012B", x"0136", x"014B", x"016F", x"018C", x"0199", x"019B", x"01A5", x"01AC", x"01B7", x"01D3", x"01D8", x"01CF", x"01BF", x"01AF", x"0198", x"0198", x"019D", x"019F", x"01A1", x"01A3", x"019F", x"018E", x"018A", x"0181", x"0175", x"017D", x"0182", x"018D", x"0187", x"0190", x"017D", x"0173", x"0163", x"014B", x"0128", x"0109", x"00E4", x"00C9", x"00C4", x"00C8", x"00D2", x"00E6", x"00EE", x"00EC", x"00EA", x"00EF", x"00FF", x"011D", x"0154", x"017D", x"019E", x"01B6", x"01C3", x"01C6", x"01CE", x"01D5", x"01C5", x"01B6", x"01A5", x"0191", x"0188", x"0192", x"019D", x"019E", x"01A2", x"019C", x"018E", x"017B", x"0170", x"015F", x"0155", x"015C", x"0160", x"0160", x"015F", x"0158", x"0144", x"0142", x"0135", x"0134", x"012A", x"0128", x"011C", x"0117", x"011D", x"0127", x"013D", x"0151", x"0166", x"0170", x"017C", x"018B", x"019A", x"01B7", x"01D9", x"01E3", x"01EE", x"01E6", x"01DB", x"01D0", x"01D2", x"01D8", x"01D9", x"01D8", x"01DC", x"01D2", x"01DD", x"01F1", x"0202", x"0215", x"0225", x"0233", x"022D", x"0233", x"022D", x"0228", x"0225", x"022F", x"0234", x"0238", x"0241", x"0235", x"0235", x"0224", x"0221", x"020A", x"01F8", x"01DE", x"01C9", x"01B8", x"01B4", x"01B5", x"01B4", x"01B5", x"01A0", x"0181", x"0160", x"0138", x"011D", x"0118", x"0119", x"011D", x"011F", x"0120", x"011B", x"011C", x"012C", x"0134", x"0134", x"0130", x"0129", x"0117", x"0121", x"0127", x"012A", x"0124", x"011B", x"0104", x"00E8", x"00D7", x"00C8", x"00BD", x"00C6", x"00D7", x"00ED", x"0101", x"0119", x"0124", x"012F", x"013D", x"0147", x"014D", x"0150", x"0151", x"0147", x"014B", x"014C", x"0157", x"015D", x"0169", x"0160", x"015B", x"0153", x"0150", x"0157", x"0171", x"0182", x"0189", x"018E", x"0183", x"0174", x"0175", x"0179", x"0178", x"0170", x"016B", x"0151", x"0140", x"0138", x"0132", x"0126", x"011B", x"010E", x"00F5", x"00E1", x"00DB", x"00CA", x"00C8", x"00CD", x"00DA", x"00DD", x"00EC", x"00EE", x"00E9", x"00E3", x"00DD", x"00CF", x"00C1", x"00B3", x"009B", x"0083", x"0075", x"0063", x"0064", x"0066", x"006E", x"006A", x"006B", x"0064", x"0067", x"0078", x"00A3", x"00C7", x"00EE", x"010F", x"011B", x"0121", x"0137", x"0144", x"0147", x"014A", x"0140", x"0135", x"0127", x"0133", x"012D", x"012A", x"0129", x"011C", x"010A", x"00FD", x"00F6", x"00E6", x"00E9", x"00E4", x"00ED", x"00E1", x"00E0", x"00CB", x"00AD", x"0092", x"0072", x"0055", x"003D", x"002C", x"0014", x"0006", x"0001", x"FFF2", x"FFFF", x"FFFD", x"0002", x"FFFE", x"FFFB", x"FFF1", x"FFF2", x"0004", x"001E", x"002E", x"0042", x"0042", x"0035", x"002D", x"002B", x"002A", x"0025", x"002B", x"0024", x"001F", x"0028", x"003C", x"0048", x"005B", x"0066", x"0065", x"005E", x"0060", x"005F", x"005C", x"0066", x"0072", x"0077", x"007D", x"007D", x"0075", x"0068", x"005E", x"0054", x"0047", x"0042", x"002F", x"0024", x"0013", x"0012", x"0009", x"000A", x"0006", x"FFF1", x"FFE0", x"FFB8", x"FFA2", x"FF8D", x"FF92", x"FF9D", x"FFAD", x"FFBA", x"FFC6", x"FFBE", x"FFCA", x"FFD1", x"FFDE", x"FFE4", x"FFED", x"FFE0", x"FFDE", x"FFE2", x"FFED", x"FFEF", x"FFF1", x"FFE9", x"FFD0", x"FFBA", x"FFA6", x"FF8D", x"FF76", x"FF6C", x"FF67", x"FF6A", x"FF75", x"FF7E", x"FF81", x"FF82", x"FF89", x"FF8D", x"FF94", x"FF9D", x"FFA3", x"FFA0", x"FFA6", x"FFAA", x"FFB4", x"FFC0", x"FFCF", x"FFD2", x"FFD6", x"FFDA", x"FFD3", x"FFDF", x"FFEF", x"FFFD", x"000E", x"0018", x"001D", x"0011", x"0016", x"0013", x"000D", x"0006", x"FFFF", x"FFE6", x"FFE3", x"FFDF", x"FFE8", x"FFE0", x"FFE5", x"FFD3", x"FFC1", x"FFB1", x"FFAE", x"FFA0", x"FFA1", x"FF9F", x"FFA7", x"FFA0", x"FFB1", x"FF9F", x"FF9A", x"FF7D", x"FF70", x"FF4F", x"FF38", x"FF23", x"FF05", x"FEEC", x"FEDB", x"FEC4", x"FEC0", x"FEB8", x"FEB5", x"FEAB", x"FEA8", x"FE9F", x"FEA0", x"FEB3", x"FECA", x"FEEC", x"FF11", x"FF2C", x"FF3B", x"FF44", x"FF51", x"FF5B", x"FF60", x"FF6C", x"FF69", x"FF5C", x"FF5E", x"FF58", x"FF4E", x"FF44", x"FF34", x"FF14", x"FEF7", x"FEDC", x"FEC8", x"FEB0", x"FEAD", x"FEA7", x"FEA8", x"FEA9", x"FEA4", x"FE97", x"FE83", x"FE76", x"FE64", x"FE5C", x"FE56", x"FE59", x"FE52", x"FE5C", x"FE5F", x"FE6A", x"FE82", x"FE94", x"FEAA", x"FEB8", x"FEC8", x"FED1", x"FEDE", x"FEF7", x"FF08", x"FF23", x"FF35", x"FF41", x"FF38", x"FF36", x"FF20", x"FF19", x"FEFF", x"FEF9", x"FEE4", x"FEDC", x"FEDF", x"FEE8", x"FEF3", x"FF03", x"FF09", x"FF0C", x"FF09", x"FF08", x"FF0A", x"FF09", x"FF19", x"FF28", x"FF37", x"FF50", x"FF55", x"FF60", x"FF50", x"FF48", x"FF2A", x"FF1D", x"FEFF", x"FEEE", x"FEDC", x"FEC9", x"FECA", x"FEC4", x"FEC4", x"FEBA", x"FEA9", x"FE8C", x"FE70", x"FE4C", x"FE40", x"FE36", x"FE3F", x"FE4E", x"FE66", x"FE73", x"FE83", x"FE8A", x"FE90", x"FE88", x"FE86", x"FE77", x"FE65", x"FE5C", x"FE56", x"FE53", x"FE51", x"FE4A", x"FE40", x"FE29", x"FE1A", x"FE11", x"FE02", x"FE0A", x"FE14", x"FE2E", x"FE46", x"FE6D", x"FE84", x"FE95", x"FE9C", x"FEA2", x"FEA5", x"FEA3", x"FEAE", x"FEA5", x"FEA6", x"FEA1", x"FEA1", x"FEA0", x"FEA3", x"FEA8", x"FEA1", x"FEA5", x"FE9D", x"FE9F", x"FE9F", x"FEAD", x"FEB8", x"FECB", x"FEDE", x"FEEC", x"FEF5", x"FEFF", x"FF01", x"FEFB", x"FEF4", x"FEE8", x"FED4", x"FEC7", x"FEC0", x"FEB5", x"FEB3", x"FEA8", x"FE9A", x"FE82", x"FE6D", x"FE5D", x"FE44", x"FE43", x"FE3C", x"FE40", x"FE47", x"FE50", x"FE58", x"FE53", x"FE58", x"FE4F", x"FE4E", x"FE49", x"FE42", x"FE31", x"FE26", x"FE11", x"FE0D", x"FE07", x"FE09", x"FE0D", x"FE0E", x"FE0F", x"FE12", x"FE19", x"FE31", x"FE4B", x"FE73", x"FEA1", x"FECD", x"FEEE", x"FF10", x"FF27", x"FF34", x"FF39", x"FF40", x"FF2F", x"FF2B", x"FF20", x"FF1D", x"FF13", x"FF0E", x"FEFC", x"FEE1", x"FEC3", x"FEB0", x"FE97", x"FE8F", x"FE8D", x"FE94", x"FE95", x"FEA7", x"FEA5", x"FEA5", x"FE93", x"FE8B", x"FE73", x"FE6D", x"FE63", x"FE60", x"FE54", x"FE52", x"FE4C", x"FE4C", x"FE4A", x"FE4B", x"FE3C", x"FE37", x"FE2A", x"FE2A", x"FE2B", x"FE32", x"FE45", x"FE4E", x"FE68", x"FE76", x"FE84", x"FE90", x"FE8F", x"FE92", x"FE90", x"FE95", x"FE9D", x"FEB1", x"FEC9", x"FEE8", x"FEFF", x"FF14", x"FF1A", x"FF0F", x"FF05", x"FEF6", x"FEED", x"FEEC", x"FEF1", x"FEF7", x"FF05", x"FF10", x"FF20", x"FF25", x"FF29", x"FF27", x"FF1F", x"FF18", x"FF0D", x"FF07", x"FEF9", x"FEF7", x"FEE6", x"FEE8", x"FED6", x"FECD", x"FEB7", x"FE9D", x"FE80", x"FE69", x"FE51", x"FE50", x"FE48", x"FE5A", x"FE6D", x"FE83", x"FE9F", x"FEB1", x"FEC5", x"FECC", x"FED6", x"FED9", x"FED9", x"FEE7", x"FEF5", x"FF0B", x"FF17", x"FF23", x"FF17", x"FF0D", x"FEF5", x"FEE6", x"FECE", x"FEC7", x"FEC1", x"FEC6", x"FED1", x"FEE9", x"FEF4", x"FF00", x"FF00", x"FEFF", x"FEF6", x"FEF6", x"FEFA", x"FEFB", x"FEFB", x"FF02", x"FF03", x"FF0C", x"FF12", x"FF23", x"FF25", x"FF2A", x"FF30", x"FF28", x"FF31", x"FF36", x"FF47", x"FF5C", x"FF75", x"FF92", x"FFA1", x"FFB3", x"FFB3", x"FFAD", x"FFA9", x"FF9B", x"FF93", x"FF8E", x"FF93", x"FF94", x"FF97", x"FF96", x"FF81", x"FF71", x"FF50", x"FF39", x"FF20", x"FF16", x"FF0C", x"FF0C", x"FF06", x"FF0F", x"FF0A", x"FF12", x"FF0D", x"FF0D", x"FF06", x"FF04", x"FF00", x"FEF6", x"FEF5", x"FEE8", x"FEE6", x"FEE4", x"FEEA", x"FEF2", x"FEF9", x"FEFF", x"FEFF", x"FF01", x"FF01", x"FF11", x"FF1A", x"FF3C", x"FF4F", x"FF6B", x"FF82", x"FF92", x"FF9C", x"FFA2", x"FFA0", x"FF9F", x"FF9B", x"FFA4", x"FFAC", x"FFBD", x"FFC8", x"FFD3", x"FFC7", x"FFC3", x"FFB1", x"FFAB", x"FFA7", x"FFAE", x"FFB3", x"FFB5", x"FFBC", x"FFBB", x"FFB3", x"FFAE", x"FF9E", x"FF90", x"FF83", x"FF7D", x"FF77", x"FF74", x"FF75", x"FF7F", x"FF8B", x"FFA1", x"FFB9", x"FFCA", x"FFDD", x"FFEB", x"FFF8", x"0009", x"0014", x"0027", x"0037", x"004E", x"005D", x"006D", x"0070", x"0067", x"005C", x"0048", x"003A", x"002B", x"002A", x"0032", x"0040", x"0057", x"0068", x"006F", x"0072", x"006E", x"006F", x"0074", x"0082", x"0093", x"00A1", x"00B8", x"00C4", x"00D4", x"00DB", x"00DD", x"00D6", x"00CE", x"00C1", x"00B7", x"00A5", x"009A", x"0089", x"0080", x"0072", x"006B", x"005D", x"004B", x"003B", x"0021", x"000E", x"FFF8", x"FFF0", x"FFEA", x"FFFF", x"0010", x"0029", x"0045", x"0053", x"0060", x"0060", x"005E", x"0050", x"0041", x"0039", x"0031", x"0036", x"003F", x"0041", x"003C", x"002C", x"001F", x"000E", x"0007", x"000A", x"0011", x"001F", x"002F", x"0048", x"0055", x"006C", x"0076", x"0075", x"007B", x"006E", x"0072", x"0067", x"0065", x"0064", x"0062", x"0066", x"0076", x"0082", x"008F", x"00A0", x"00A2", x"00B1", x"00B8", x"00C5", x"00DE", x"00F1", x"0113", x"012A", x"0143", x"0150", x"0154", x"014D", x"0141", x"0129", x"011B", x"010D", x"0106", x"0102", x"00FE", x"00F4", x"00DB", x"00C5", x"00A2", x"008A", x"007C", x"0075", x"007F", x"008A", x"009E", x"00AB", x"00C4", x"00D9", x"00F0", x"00FC", x"0108", x"0103", x"00FD", x"00ED", x"00DF", x"00CE", x"00C3", x"00B7", x"00B2", x"00AF", x"00AC", x"00AE", x"00AA", x"00B1", x"00BC", x"00C8", x"00E7", x"010E", x"0132", x"0163", x"0189", x"01AE", x"01BE", x"01CD", x"01C2", x"01BD", x"01AF", x"01AE", x"01A7", x"01A9", x"01A7", x"019C", x"0185", x"0174", x"015A", x"014C", x"0143", x"0141", x"0144", x"0142", x"014D", x"0148", x"0150", x"014A", x"0147", x"0138", x"012F", x"0127", x"0116", x"010F", x"00FD", x"00F8", x"00E8", x"00F0", x"00EC", x"00EF", x"00F3", x"00E7", x"00EE", x"00EA", x"00EE", x"00FA", x"0102", x"0114", x"0121", x"0131", x"013B", x"0142", x"0144", x"0142", x"0144", x"0143", x"0154", x"0160", x"017B", x"0187", x"0197", x"0195", x"018D", x"0183", x"0177", x"016D", x"016D", x"016B", x"016E", x"017E", x"0185", x"019A", x"01A9", x"01BC", x"01C5", x"01CE", x"01CF", x"01CE", x"01C1", x"01B9", x"01A5", x"018F", x"0182", x"0170", x"015F", x"0151", x"013D", x"0125", x"0109", x"00F5", x"00DF", x"00DA", x"00E2", x"00EF", x"0108", x"011B", x"013C", x"014D", x"016A", x"017A", x"0181", x"0181", x"0186", x"018D", x"0194", x"01A1", x"01A5", x"0197", x"018C", x"016F", x"015B", x"013B", x"0137", x"0122", x"0123", x"0120", x"012B", x"012A", x"0137", x"013D", x"0140", x"0149", x"0151", x"015E", x"0168", x"0174", x"0184", x"0192", x"01A9", x"01BF", x"01CF", x"01D7", x"01E0", x"01D6", x"01D8", x"01D4", x"01D2", x"01D9", x"01E3", x"01F2", x"01FD", x"020E", x"0217", x"021E", x"0220", x"021F", x"0216", x"0212", x"020C", x"0209", x"0205", x"0207", x"01F7", x"01E7", x"01CA", x"01B4", x"0193", x"0189", x"0178", x"0170", x"016A", x"016C", x"0169", x"016B", x"0170", x"0170", x"016D", x"016D", x"0169", x"0163", x"0155", x"0146", x"012E", x"011E", x"010F", x"0108", x"00FC", x"00FD", x"00F0", x"00EB", x"00E2", x"00E4", x"00E4", x"00F2", x"0107", x"0118", x"0130", x"014E", x"0160", x"017B", x"0184", x"018A", x"0181", x"017A", x"0177", x"0176", x"0172", x"0178", x"0167", x"0158", x"0145", x"012A", x"0117", x"0100", x"00F8", x"00E1", x"00DC", x"00D5", x"00CE", x"00CA", x"00C4", x"00BA", x"00B0", x"00A6", x"00A4", x"0098", x"009E", x"0093", x"0099", x"009E", x"00AF", x"00BC", x"00D3", x"00D8", x"00E9", x"00DE", x"00E8", x"00DD", x"00EA", x"00EA", x"00F9", x"00F8", x"0100", x"00FE", x"00F8", x"00FA", x"00F2", x"00ED", x"00E4", x"00E4", x"00E1", x"00EE", x"00F8", x"010B", x"010E", x"0114", x"0110", x"010F", x"010D", x"0119", x"011E", x"0128", x"0135", x"013D", x"014A", x"014F", x"015B", x"014E", x"014B", x"0136", x"0124", x"0108", x"00F8", x"00D5", x"00C2", x"00A8", x"009D", x"0087", x"007A", x"0068", x"0051", x"003D", x"002A", x"001C", x"0014", x"001E", x"0021", x"0031", x"003A", x"004B", x"0054", x"005B", x"005C", x"004F", x"0042", x"0035", x"002D", x"0029", x"0032", x"0031", x"002F", x"0028", x"0020", x"000C", x"0009", x"FFFE", x"0001", x"0000", x"0015", x"001D", x"0034", x"0040", x"004F", x"0051", x"0059", x"0054", x"0051", x"0047", x"0043", x"0037", x"002F", x"0029", x"0026", x"0025", x"002A", x"002D", x"0031", x"0035", x"0037", x"0039", x"0048", x"0056", x"006A", x"0076", x"008B", x"008C", x"0095", x"0098", x"0095", x"008A", x"0081", x"0070", x"005F", x"0054", x"0047", x"0035", x"0011", x"FFF6", x"FFC9", x"FFA8", x"FF8C", x"FF73", x"FF5B", x"FF51", x"FF51", x"FF58", x"FF6C", x"FF83", x"FF93", x"FF9C", x"FFA6", x"FFAD", x"FFB0", x"FFAC", x"FFA7", x"FF90", x"FF88", x"FF7B", x"FF7D", x"FF7C", x"FF80", x"FF82", x"FF7D", x"FF81", x"FF7E", x"FF84", x"FF95", x"FFAA", x"FFC9", x"FFE7", x"0008", x"0020", x"0038", x"0049", x"0051", x"0049", x"0041", x"002A", x"0018", x"000D", x"0001", x"FFF1", x"FFE0", x"FFC5", x"FFA5", x"FF8A", x"FF74", x"FF66", x"FF59", x"FF5D", x"FF5E", x"FF61", x"FF68", x"FF65", x"FF63", x"FF54", x"FF56", x"FF45", x"FF40", x"FF34", x"FF22", x"FF12", x"FF06", x"FEF7", x"FEED", x"FEE5", x"FEDF", x"FED3", x"FECC", x"FEC0", x"FEB5", x"FEBC", x"FEC1", x"FED2", x"FEDA", x"FEE6", x"FEEB", x"FEEC", x"FEF7", x"FF09", x"FF0F", x"FF21", x"FF2E", x"FF35", x"FF45", x"FF59", x"FF62", x"FF68", x"FF65", x"FF5C", x"FF4E", x"FF3E", x"FF3C", x"FF2B", x"FF2A", x"FF31", x"FF3A", x"FF4D", x"FF62", x"FF72", x"FF7A", x"FF80", x"FF88", x"FF83", x"FF80", x"FF6F", x"FF56", x"FF39", x"FF22", x"FF09", x"FEF6", x"FEE3", x"FECD", x"FEB3", x"FE95", x"FE7D", x"FE61", x"FE54", x"FE4B", x"FE4E", x"FE52", x"FE68", x"FE75", x"FE8E", x"FEA8", x"FEB6", x"FEC6", x"FECB", x"FED1", x"FECB", x"FED4", x"FEDD", x"FEDD", x"FEE1", x"FEDB", x"FEC3", x"FEB0", x"FE9A", x"FE87", x"FE79", x"FE73", x"FE7B", x"FE83", x"FE8F", x"FEA1", x"FE9F", x"FEA0", x"FEA0", x"FE9A", x"FE98", x"FE9F", x"FE9A", x"FE9F", x"FE9B", x"FEA4", x"FEAD", x"FEBE", x"FECF", x"FEDB", x"FEE0", x"FEE0", x"FEDF", x"FEDC", x"FEF0", x"FEFD", x"FF10", x"FF1E", x"FF2C", x"FF2C", x"FF3B", x"FF44", x"FF49", x"FF46", x"FF47", x"FF37", x"FF29", x"FF25", x"FF19", x"FF08", x"FEF1", x"FED3", x"FEA8", x"FE82", x"FE5C", x"FE41", x"FE1B", x"FE18", x"FE0B", x"FE14", x"FE24", x"FE34", x"FE49", x"FE54", x"FE6D", x"FE7B", x"FE83", x"FE85", x"FE77", x"FE5F", x"FE4D", x"FE38", x"FE30", x"FE28", x"FE26", x"FE22", x"FE1D", x"FE16", x"FE0A", x"FE07", x"FDFF", x"FE06", x"FE0E", x"FE24", x"FE30", x"FE41", x"FE59", x"FE60", x"FE73", x"FE79", x"FE7F", x"FE76", x"FE72", x"FE7E", x"FE7E", x"FE93", x"FE93", x"FE99", x"FE82", x"FE80", x"FE70", x"FE5E", x"FE53", x"FE49", x"FE47", x"FE4A", x"FE55", x"FE5C", x"FE59", x"FE57", x"FE58", x"FE4A", x"FE51", x"FE43", x"FE3D", x"FE2D", x"FE2F", x"FE2F", x"FE40", x"FE51", x"FE65", x"FE72", x"FE7E", x"FE80", x"FE80", x"FE83", x"FE88", x"FE8E", x"FE95", x"FE9E", x"FE9B", x"FE9E", x"FE9D", x"FEA0", x"FEA5", x"FEAA", x"FEB4", x"FEB1", x"FEC0", x"FECD", x"FED2", x"FEDE", x"FEDE", x"FEDA", x"FED7", x"FED2", x"FED3", x"FECB", x"FECF", x"FEDC", x"FEEA", x"FF06", x"FF1C", x"FF34", x"FF33", x"FF42", x"FF40", x"FF3E", x"FF38", x"FF23", x"FF08", x"FEE4", x"FEC2", x"FEA7", x"FE8B", x"FE7C", x"FE67", x"FE59", x"FE42", x"FE32", x"FE1D", x"FE1F", x"FE18", x"FE2C", x"FE39", x"FE51", x"FE60", x"FE77", x"FE95", x"FEA5", x"FEC0", x"FECB", x"FEC6", x"FEC2", x"FEBB", x"FEC2", x"FEBD", x"FEC8", x"FEC1", x"FEAD", x"FE9B", x"FE8B", x"FE78", x"FE62", x"FE62", x"FE5C", x"FE62", x"FE75", x"FE87", x"FE91", x"FE9E", x"FEA9", x"FEB1", x"FEBB", x"FEC4", x"FEC3", x"FEBB", x"FEB2", x"FEB4", x"FEB2", x"FEC7", x"FED8", x"FEE7", x"FEF2", x"FEF1", x"FEF3", x"FEF0", x"FEFB", x"FF06", x"FF1A", x"FF2B", x"FF3A", x"FF42", x"FF49", x"FF4D", x"FF49", x"FF49", x"FF3B", x"FF25", x"FF0D", x"FEFC", x"FEE6", x"FED4", x"FEC2", x"FEA3", x"FE80", x"FE5D", x"FE44", x"FE25", x"FE1E", x"FE20", x"FE28", x"FE49", x"FE67", x"FE96", x"FEAF", x"FED6", x"FEEA", x"FEFB", x"FF08", x"FF0A", x"FF0A", x"FEF9", x"FEF4", x"FEEC", x"FEEE", x"FEF8", x"FEFF", x"FF05", x"FF05", x"FF01", x"FEF7", x"FEF7", x"FEF1", x"FF01", x"FF0F", x"FF31", x"FF46", x"FF63", x"FF80", x"FF91", x"FFAA", x"FFBB", x"FFC2", x"FFBB", x"FFBE", x"FFB4", x"FFB0", x"FFAF", x"FFA4", x"FF95", x"FF7A", x"FF69", x"FF53", x"FF3A", x"FF2A", x"FF1E", x"FF0D", x"FF11", x"FF1B", x"FF1E", x"FF24", x"FF25", x"FF26", x"FF26", x"FF28", x"FF25", x"FF16", x"FF03", x"FEF0", x"FEEA", x"FEE6", x"FEF3", x"FEFA", x"FF00", x"FF04", x"FF07", x"FF02", x"FF04", x"FF07", x"FF0F", x"FF1D", x"FF2E", x"FF33", x"FF43", x"FF4D", x"FF61", x"FF78", x"FF93", x"FFA1", x"FFB3", x"FFBF", x"FFD5", x"FFE3", x"FFFD", x"000F", x"000A", x"0013", x"0007", x"0000", x"FFEF", x"FFEA", x"FFE3", x"FFE5", x"FFF9", x"0012", x"0029", x"003A", x"0051", x"0055", x"0060", x"005F", x"0055", x"003A", x"001F", x"0005", x"FFE5", x"FFE8", x"FFDD", x"FFE0", x"FFD3", x"FFCA", x"FFB5", x"FFA3", x"FF99", x"FF91", x"FF98", x"FF9E", x"FFAF", x"FFB6", x"FFCB", x"FFDF", x"FFF2", x"0009", x"001A", x"0022", x"0022", x"0028", x"0028", x"0024", x"002B", x"001A", x"0009", x"FFF0", x"FFD9", x"FFC0", x"FFAE", x"FFAB", x"FFA6", x"FFAC", x"FFC8", x"FFDC", x"FFF2", x"0008", x"001E", x"002C", x"0040", x"0059", x"005F", x"0068", x"0069", x"0069", x"0070", x"007C", x"0096", x"00A3", x"00B5", x"00BF", x"00C3", x"00CA", x"00D7", x"00E1", x"00F1", x"00FE", x"010C", x"010A", x"011E", x"011B", x"0125", x"012A", x"012B", x"0125", x"0119", x"0116", x"0103", x"00F7", x"00EA", x"00CC", x"00B3", x"009D", x"0081", x"0068", x"0055", x"0046", x"003C", x"0041", x"0056", x"006A", x"0080", x"009A", x"00AB", x"00B5", x"00BE", x"00C0", x"00AA", x"0093", x"0076", x"0057", x"0048", x"0043", x"0047", x"004B", x"004B", x"0049", x"003B", x"003F", x"0037", x"0045", x"0055", x"006B", x"0081", x"009B", x"00AD", x"00C7", x"00D4", x"00E7", x"00EE", x"00EA", x"00EC", x"00E7", x"00E2", x"00E8", x"00E3", x"00E4", x"00D3", x"00D4", x"00BD", x"00B4", x"00A8", x"00A4", x"009B", x"00AC", x"00B1", x"00C5", x"00C4", x"00D1", x"00C9", x"00C8", x"00C7", x"00BE", x"00B1", x"00A1", x"0098", x"008C", x"0099", x"00AC", x"00C6", x"00D6", x"00E4", x"00E1", x"00DC", x"00DE", x"00DF", x"00E5", x"00F6", x"00F6", x"0102", x"0107", x"011A", x"0129", x"0143", x"0158", x"016E", x"0173", x"0182", x"0187", x"0186", x"018D", x"018B", x"017D", x"017B", x"016E", x"0164", x"0154", x"014E", x"0145", x"0145", x"0158", x"0163", x"0176", x"017E", x"0189", x"0192", x"0191", x"0197", x"0188", x"0171", x"0155", x"0138", x"0121", x"0113", x"011C", x"0115", x"011E", x"0117", x"010A", x"00FD", x"00F3", x"00EC", x"00F0", x"00F6", x"0103", x"010F", x"0123", x"013A", x"014D", x"016A", x"0176", x"017E", x"0178", x"0176", x"016D", x"0169", x"0168", x"0160", x"0156", x"014A", x"0144", x"012A", x"0122", x"010D", x"0102", x"00FB", x"0105", x"010E", x"011A", x"0131", x"0134", x"0141", x"0147", x"0150", x"014E", x"0142", x"0133", x"0121", x"0114", x"011F", x"0125", x"0137", x"0144", x"0144", x"0145", x"013A", x"0146", x"0148", x"015B", x"0170", x"0184", x"0193", x"01AF", x"01BB", x"01D1", x"01E0", x"01E9", x"01E0", x"01DC", x"01C8", x"01B2", x"0194", x"017C", x"014C", x"012F", x"0107", x"00E1", x"00C1", x"00A5", x"009A", x"0093", x"00A1", x"00BE", x"00D8", x"00FC", x"0119", x"0136", x"014E", x"0167", x"0173", x"0172", x"0169", x"0156", x"0145", x"013D", x"013F", x"0148", x"0151", x"0156", x"0154", x"0149", x"013E", x"0132", x"0136", x"013D", x"014A", x"0154", x"0161", x"016F", x"017C", x"019D", x"01B0", x"01C5", x"01C9", x"01CC", x"01C0", x"01BA", x"01B5", x"01AE", x"01A1", x"0199", x"0188", x"0175", x"0163", x"0154", x"013B", x"012E", x"0123", x"011E", x"011C", x"0122", x"0127", x"0126", x"012E", x"012F", x"012A", x"011A", x"0109", x"00EA", x"00D7", x"00CB", x"00CA", x"00D5", x"00DA", x"00E3", x"00DC", x"00DA", x"00DA", x"00D8", x"00E5", x"00F1", x"00FE", x"0109", x"0117", x"0126", x"0133", x"014E", x"015C", x"016C", x"0173", x"0178", x"0180", x"0181", x"0190", x"018D", x"018C", x"0186", x"017A", x"0167", x"0157", x"014A", x"0139", x"013B", x"013D", x"0152", x"015D", x"017A", x"0183", x"0192", x"0195", x"0194", x"0185", x"0170", x"0153", x"012F", x"0116", x"00FA", x"00EE", x"00DD", x"00D6", x"00C2", x"00AC", x"0094", x"0079", x"0065", x"0059", x"0056", x"0058", x"005B", x"0066", x"0070", x"0084", x"00A1", x"00B8", x"00CF", x"00DD", x"00E2", x"00E1", x"00DE", x"00D8", x"00CD", x"00C1", x"00B7", x"00A3", x"0098", x"0082", x"007A", x"0065", x"006B", x"0064", x"006E", x"0074", x"0088", x"008C", x"009B", x"00A6", x"00B3", x"00B8", x"00BE", x"00B4", x"00A6", x"009D", x"00A3", x"00AC", x"00C8", x"00D9", x"00ED", x"00ED", x"00FA", x"00F7", x"0103", x"0107", x"0116", x"0118", x"011D", x"0120", x"0123", x"0124", x"0128", x"011F", x"011A", x"0102", x"00E9", x"00CC", x"00AE", x"009C", x"0080", x"0073", x"0056", x"003E", x"001F", x"000B", x"FFF1", x"FFF6", x"FFF2", x"0004", x"0013", x"002A", x"0044", x"005A", x"0072", x"0082", x"0088", x"0080", x"006D", x"0049", x"0027", x"000A", x"FFF3", x"FFE9", x"FFE2", x"FFD2", x"FFC1", x"FFAA", x"FF98", x"FF8D", x"FF87", x"FF93", x"FF98", x"FFA9", x"FFB5", x"FFC4", x"FFD7", x"FFF2", x"000D", x"0027", x"003A", x"003C", x"003E", x"0035", x"0036", x"002C", x"002B", x"001F", x"0017", x"0008", x"FFFE", x"FFF8", x"FFF2", x"FFF4", x"FFF9", x"FFF9", x"0000", x"0005", x"0008", x"000D", x"0010", x"0011", x"0008", x"FFFE", x"FFE7", x"FFCF", x"FFB7", x"FFA9", x"FF9E", x"FFA2", x"FFA0", x"FFAB", x"FFA3", x"FFA9", x"FF9B", x"FF9A", x"FF92", x"FF91", x"FF8F", x"FF8D", x"FF94", x"FF98", x"FFA7", x"FFB9", x"FFCE", x"FFE2", x"FFF4", x"0000", x"0004", x"0003", x"0003", x"0002", x"0002", x"0002", x"FFFD", x"FFF4", x"FFE6", x"FFDC", x"FFD4", x"FFD5", x"FFDA", x"FFE5", x"FFF4", x"0003", x"0012", x"0020", x"0021", x"0025", x"0016", x"0003", x"FFDF", x"FFBB", x"FF93", x"FF78", x"FF5B", x"FF53", x"FF41", x"FF3A", x"FF2B", x"FF1B", x"FF0F", x"FF03", x"FF05", x"FF09", x"FF19", x"FF28", x"FF3F", x"FF4F", x"FF65", x"FF78", x"FF8A", x"FF95", x"FF97", x"FF96", x"FF81", x"FF73", x"FF5C", x"FF4B", x"FF42", x"FF31", x"FF24", x"FF09", x"FEF1", x"FEDB", x"FECF", x"FEC5", x"FECC", x"FECD", x"FED9", x"FEE2", x"FEF3", x"FF02", x"FF17", x"FF27", x"FF32", x"FF37", x"FF2F", x"FF25", x"FF16", x"FF0D", x"FF0E", x"FF18", x"FF1D", x"FF2A", x"FF25", x"FF2B", x"FF28", x"FF2C", x"FF33", x"FF37", x"FF3F", x"FF43", x"FF4C", x"FF55", x"FF5B", x"FF6C", x"FF6B", x"FF6E", x"FF66", x"FF53", x"FF3C", x"FF1C", x"FEFB", x"FEE3", x"FEBF", x"FEA7", x"FE83", x"FE66", x"FE4B", x"FE41", x"FE41", x"FE4D", x"FE5F", x"FE77", x"FE96", x"FEB4", x"FEDB", x"FEF9", x"FF13", x"FF26", x"FF2F", x"FF28", x"FF1B", x"FF06", x"FEF2", x"FEE3", x"FEDF", x"FEDB", x"FEDB", x"FED6", x"FECF", x"FEC2", x"FEB8", x"FEB0", x"FEAE", x"FEB5", x"FEBB", x"FECC", x"FEDC", x"FEF3", x"FF08", x"FF22", x"FF33", x"FF46", x"FF48", x"FF47", x"FF3E", x"FF33", x"FF23", x"FF15", x"FF09", x"FEF7", x"FEE4", x"FEC9", x"FEB5", x"FE99", x"FE8E", x"FE7C", x"FE7C", x"FE79", x"FE7B", x"FE83", x"FE8F", x"FE9A", x"FEAB", x"FEAF", x"FEB3", x"FEAA", x"FE98", x"FE88", x"FE6A", x"FE61", x"FE54", x"FE4D", x"FE4E", x"FE4E", x"FE4C", x"FE4E", x"FE4C", x"FE53", x"FE60", x"FE6C", x"FE81", x"FE91", x"FEA7", x"FEBD", x"FED5", x"FEEF", x"FF05", x"FF17", x"FF25", x"FF31", x"FF38", x"FF38", x"FF39", x"FF33", x"FF29", x"FF20", x"FF05", x"FEF0", x"FED5", x"FEC5", x"FEB9", x"FEBA", x"FEBE", x"FEC1", x"FEC8", x"FED5", x"FEE3", x"FEF2", x"FF00", x"FF04", x"FEFE", x"FEEA", x"FEDB", x"FEBD", x"FEB0", x"FEA0", x"FE9B", x"FE95", x"FE8C", x"FE86", x"FE71", x"FE66", x"FE51", x"FE4F", x"FE3F", x"FE47", x"FE3F", x"FE48", x"FE52", x"FE66", x"FE78", x"FE93", x"FE9B", x"FEAC", x"FEAA", x"FEAB", x"FEA3", x"FE9A", x"FE8C", x"FE83", x"FE75", x"FE6A", x"FE55", x"FE4B", x"FE3C", x"FE3A", x"FE3B", x"FE44", x"FE51", x"FE5A", x"FE70", x"FE81", x"FEA0", x"FEBA", x"FED8", x"FEEF", x"FEFD", x"FF04", x"FF02", x"FEFE", x"FEFA", x"FEFB", x"FF04", x"FF0E", x"FF1E", x"FF2A", x"FF31", x"FF3B", x"FF3E", x"FF47", x"FF4D", x"FF51", x"FF5B", x"FF5A", x"FF66", x"FF62", x"FF69", x"FF61", x"FF60", x"FF59", x"FF4D", x"FF45", x"FF33", x"FF24", x"FF13", x"FEFB", x"FEEE", x"FED3", x"FEC1", x"FEAD", x"FEA2", x"FE99", x"FE9F", x"FE9D", x"FEAE", x"FEB8", x"FED4", x"FEE6", x"FF06", x"FF13", x"FF30", x"FF31", x"FF3D", x"FF28", x"FF24", x"FEFF", x"FEF5", x"FEDC", x"FED3", x"FEC6", x"FEB8", x"FEB0", x"FE98", x"FE8C", x"FE81", x"FE7D", x"FE80", x"FE86", x"FE92", x"FEA0", x"FEB3", x"FECE", x"FEE3", x"FEFD", x"FF15", x"FF27", x"FF31", x"FF3C", x"FF3B", x"FF3D", x"FF3A", x"FF32", x"FF28", x"FF1A", x"FF0D", x"FF04", x"FEF4", x"FEF8", x"FEEF", x"FEF4", x"FEF4", x"FEF1", x"FEF6", x"FEEF", x"FEF6", x"FEF7", x"FEFC", x"FEFA", x"FEEA", x"FEDB", x"FEBF", x"FEB1", x"FE9E", x"FEA4", x"FEA1", x"FEB4", x"FEBC", x"FEC8", x"FECB", x"FED2", x"FEDA", x"FEE1", x"FEF4", x"FEFF", x"FF0C", x"FF18", x"FF28", x"FF3F", x"FF54", x"FF75", x"FF83", x"FF99", x"FF9E", x"FFAB", x"FFAE", x"FFAD", x"FFAC", x"FF9F", x"FF91", x"FF84", x"FF6E", x"FF68", x"FF59", x"FF60", x"FF60", x"FF6A", x"FF72", x"FF7F", x"FF8C", x"FF9E", x"FFAE", x"FFC4", x"FFCB", x"FFCA", x"FFBD", x"FFA5", x"FF91", x"FF79", x"FF68", x"FF5A", x"FF4C", x"FF46", x"FF3B", x"FF31", x"FF2D", x"FF23", x"FF2B", x"FF31", x"FF46", x"FF58", x"FF6C", x"FF83", x"FF9E", x"FFB5", x"FFC9", x"FFD9", x"FFE0", x"FFE2", x"FFE2", x"FFDE", x"FFDB", x"FFCC", x"FFC3", x"FFB0", x"FF9D", x"FF91", x"FF81", x"FF80", x"FF70", x"FF78", x"FF6C", x"FF6D", x"FF6D", x"FF6D", x"FF79", x"FF7E", x"FF93", x"FF9B", x"FFA4", x"FFAA", x"FFA2", x"FFA1", x"FF92", x"FF94", x"FF88", x"FF8E", x"FF91", x"FF99", x"FFAD", x"FFB1", x"FFC7", x"FFCC", x"FFDD", x"FFE6", x"FFF4", x"0002", x"000F", x"0021", x"002E", x"003C", x"003E", x"0047", x"003C", x"0036", x"0027", x"001E", x"FFFE", x"FFE7", x"FFC5", x"FFA1", x"FF82", x"FF73", x"FF60", x"FF62", x"FF62", x"FF72", x"FF7B", x"FF9C", x"FFB3", x"FFDA", x"FFFD", x"0020", x"0043", x"005C", x"0071", x"0078", x"0074", x"0068", x"005A", x"0051", x"0041", x"0046", x"0034", x"0033", x"0024", x"0014", x"000C", x"0001", x"0003", x"000B", x"0020", x"0030", x"0047", x"005F", x"007B", x"0098", x"00B4", x"00CB", x"00DD", x"00E2", x"00EC", x"00E6", x"00EA", x"00E2", x"00D5", x"00C0", x"00A5", x"0090", x"0072", x"005F", x"004A", x"003B", x"0028", x"0021", x"0016", x"0014", x"0012", x"001B", x"0021", x"0030", x"0038", x"0038", x"002E", x"0021", x"000C", x"0003", x"FFF1", x"FFF3", x"FFEC", x"FFEF", x"FFF1", x"FFF8", x"0003", x"0012", x"0026", x"0041", x"005D", x"0075", x"0094", x"00AA", x"00C7", x"00DE", x"00FE", x"010E", x"011F", x"012D", x"0134", x"013A", x"0139", x"0130", x"0123", x"0106", x"00F8", x"00E0", x"00D0", x"00C8", x"00BE", x"00B8", x"00B5", x"00B4", x"00BB", x"00C5", x"00D2", x"00E8", x"00F1", x"00FC", x"00F6", x"00EA", x"00CD", x"00BD", x"00A1", x"0094", x"007C", x"006A", x"0059", x"0045", x"003E", x"0032", x"0028", x"0026", x"0022", x"002C", x"0032", x"0042", x"0054", x"0066", x"007E", x"0097", x"00AB", x"00BD", x"00C8", x"00D3", x"00D8", x"00DB", x"00DB", x"00CF", x"00C0", x"00A8", x"009A", x"0088", x"007F", x"007A", x"007C", x"0080", x"0088", x"0093", x"00A1", x"00B4", x"00C8", x"00EA", x"00FF", x"0126", x"0133", x"0142", x"0145", x"0147", x"0146", x"014C", x"014A", x"0151", x"0153", x"0154", x"015C", x"015D", x"016A", x"016E", x"017F", x"0183", x"0183", x"0184", x"0175", x"017A", x"0162", x"0168", x"0154", x"0144", x"0139", x"0122", x"011A", x"010C", x"00FE", x"00F3", x"00DA", x"00C9", x"00BD", x"00AF", x"00B2", x"00B7", x"00BD", x"00C6", x"00D6", x"00E3", x"00F3", x"010B", x"011D", x"0137", x"0143", x"014D", x"014F", x"0141", x"013C", x"0122", x"0114", x"00FF", x"00EB", x"00D5", x"00BE", x"00AA", x"0090", x"0084", x"0074", x"0070", x"0070", x"0075", x"0077", x"0085", x"0091", x"00A8", x"00BB", x"00DF", x"00F0", x"010C", x"011C", x"0136", x"0141", x"0154", x"0156", x"014C", x"0141", x"012E", x"0124", x"0116", x"011A", x"0117", x"0120", x"011C", x"0128", x"0123", x"012C", x"012F", x"0137", x"0135", x"013B", x"0131", x"012F", x"011B", x"0113", x"0101", x"00F5", x"00E7", x"00DF", x"00D7", x"00D9", x"00DB", x"00E2", x"00EA", x"00F0", x"00F9", x"0105", x"010F", x"0119", x"0126", x"012D", x"013A", x"014B", x"015C", x"016E", x"017F", x"018C", x"0198", x"019F", x"01A4", x"01A9", x"0198", x"0191", x"017E", x"016F", x"0162", x"015C", x"0158", x"0157", x"0157", x"0159", x"015A", x"0158", x"015C", x"015E", x"015F", x"0166", x"015C", x"0159", x"0141", x"0138", x"0127", x"011C", x"0111", x"0104", x"00F7", x"00E9", x"00DF", x"00D9", x"00DA", x"00E0", x"00EF", x"0105", x"0111", x"0126", x"012D", x"013C", x"0141", x"0156", x"0159", x"0162", x"015F", x"015F", x"0159", x"0155", x"0152", x"0145", x"0130", x"0119", x"0105", x"00F2", x"00EA", x"00E8", x"00ED", x"00ED", x"00FF", x"00FC", x"0108", x"0103", x"0110", x"0114", x"011D", x"012D", x"0131", x"0136", x"0135", x"0133", x"0131", x"0125", x"0121", x"010E", x"0107", x"00FB", x"00FA", x"00F9", x"00FB", x"00FC", x"0103", x"0108", x"0107", x"0109", x"0102", x"00FF", x"00F8", x"00F9", x"00EF", x"00DE", x"00D2", x"00C2", x"00B4", x"00A9", x"00A0", x"0084", x"006A", x"0051", x"003C", x"002F", x"0036", x"003D", x"004A", x"005C", x"0073", x"0086", x"00A7", x"00BC", x"00E0", x"00EB", x"0104", x"010D", x"010B", x"010D", x"0106", x"00FB", x"00F5", x"00E3", x"00D5", x"00BB", x"00AB", x"008D", x"0080", x"006C", x"0068", x"0061", x"006D", x"0073", x"0081", x"0089", x"0096", x"009B", x"00AA", x"00BA", x"00BC", x"00C3", x"00C3", x"00C6", x"00C1", x"00D0", x"00C5", x"00BF", x"00A2", x"008C", x"006B", x"0050", x"0044", x"0033", x"002B", x"0024", x"0021", x"0015", x"0010", x"000E", x"0007", x"000C", x"000D", x"001B", x"0014", x"001E", x"0012", x"000F", x"0006", x"FFF8", x"FFEC", x"FFDF", x"FFD0", x"FFD0", x"FFCD", x"FFD7", x"FFE4", x"0002", x"0019", x"003A", x"0053", x"006B", x"007B", x"0088", x"00A0", x"00AC", x"00BB", x"00C7", x"00CE", x"00CB", x"00D5", x"00D3", x"00CD", x"00B6", x"009B", x"007B", x"0057", x"0041", x"0031", x"0020", x"0013", x"0013", x"000F", x"0011", x"0018", x"001B", x"0020", x"001E", x"0023", x"001C", x"0013", x"0008", x"FFFF", x"FFEF", x"FFEB", x"FFDB", x"FFD6", x"FFBD", x"FFB5", x"FFA0", x"FF99", x"FF85", x"FF84", x"FF7D", x"FF7D", x"FF7E", x"FF7F", x"FF7E", x"FF7B", x"FF82", x"FF88", x"FF90", x"FF96", x"FF98", x"FF9E", x"FF9A", x"FFA7", x"FFAB", x"FFA8", x"FF95", x"FF85", x"FF66", x"FF55", x"FF4F", x"FF46", x"FF4C", x"FF4B", x"FF5D", x"FF64", x"FF76", x"FF81", x"FF94", x"FF9E", x"FFB5", x"FFC8", x"FFD9", x"FFE3", x"FFF2", x"FFF8", x"FFFF", x"0003", x"0007", x"FFFF", x"FFF6", x"FFE9", x"FFDB", x"FFD3", x"FFCE", x"FFC9", x"FFD6", x"FFD0", x"FFDC", x"FFD5", x"FFD3", x"FFC1", x"FFC1", x"FFB5", x"FFAF", x"FF9E", x"FF92", x"FF7C", x"FF6E", x"FF6A", x"FF64", x"FF53", x"FF42", x"FF29", x"FF0A", x"FEFC", x"FEF6", x"FEF5", x"FEF9", x"FF07", x"FF0E", x"FF21", x"FF28", x"FF40", x"FF47", x"FF50", x"FF5E", x"FF64", x"FF65", x"FF6B", x"FF61", x"FF5E", x"FF54", x"FF4B", x"FF39", x"FF21", x"FF07", x"FEE8", x"FEC9", x"FEB1", x"FE9D", x"FE90", x"FE8C", x"FE8C", x"FE90", x"FE97", x"FEA0", x"FEA8", x"FEC2", x"FED7", x"FEF0", x"FF08", x"FF18", x"FF20", x"FF2F", x"FF3D", x"FF3C", x"FF38", x"FF2B", x"FF0F", x"FEF6", x"FEE0", x"FED2", x"FEC8", x"FEBC", x"FEB7", x"FEA8", x"FE9F", x"FE9C", x"FE92", x"FE90", x"FE84", x"FE87", x"FE7A", x"FE7F", x"FE7F", x"FE7C", x"FE7F", x"FE78", x"FE7A", x"FE70", x"FE70", x"FE64", x"FE68", x"FE60", x"FE69", x"FE69", x"FE7E", x"FE8E", x"FEA5", x"FEBF", x"FED2", x"FEDE", x"FEED", x"FEF9", x"FEFD", x"FF0B", x"FF0F", x"FF0B", x"FF0A", x"FF0A", x"FF0E", x"FF0C", x"FF0A", x"FEFD", x"FEE8", x"FED1", x"FEC5", x"FEB7", x"FEB5", x"FEB4", x"FEB9", x"FEB6", x"FEBA", x"FEBE", x"FEBA", x"FEBE", x"FEB8", x"FEB7", x"FEB0", x"FEAD", x"FEAF", x"FEA9", x"FEAF", x"FEA9", x"FEAB", x"FEA0", x"FE97", x"FE83", x"FE78", x"FE66", x"FE63", x"FE62", x"FE73", x"FE7B", x"FE95", x"FEA4", x"FEAC", x"FEB5", x"FEB6", x"FEC0", x"FEC7", x"FECF", x"FED4", x"FECD", x"FECD", x"FECB", x"FECF", x"FEC7", x"FECB", x"FEBA", x"FEA8", x"FE96", x"FE8F", x"FE84", x"FE86", x"FE81", x"FE7C", x"FE72", x"FE6A", x"FE63", x"FE58", x"FE59", x"FE53", x"FE55", x"FE54", x"FE61", x"FE63", x"FE6D", x"FE72", x"FE76", x"FE77", x"FE79", x"FE75", x"FE70", x"FE6C", x"FE6B", x"FE62", x"FE6C", x"FE72", x"FE7B", x"FE88", x"FE8A", x"FE8F", x"FE87", x"FE8D", x"FE88", x"FE88", x"FE7F", x"FE7A", x"FE61", x"FE5F", x"FE57", x"FE5A", x"FE50", x"FE4F", x"FE3D", x"FE2D", x"FE25", x"FE24", x"FE29", x"FE3B", x"FE50", x"FE62", x"FE7D", x"FE90", x"FEAD", x"FEBC", x"FED1", x"FED7", x"FED9", x"FED5", x"FED5", x"FED1", x"FED1", x"FED1", x"FEC8", x"FEBE", x"FEB0", x"FE96", x"FE84", x"FE6B", x"FE5E", x"FE50", x"FE56", x"FE63", x"FE72", x"FE8F", x"FE9D", x"FEB0", x"FEBD", x"FED6", x"FEE8", x"FEFC", x"FF11", x"FF0E", x"FF12", x"FF14", x"FF13", x"FF19", x"FF13", x"FF08", x"FEE8", x"FECD", x"FEB2", x"FEA1", x"FE96", x"FE94", x"FE98", x"FE90", x"FE93", x"FE94", x"FE8D", x"FE95", x"FE97", x"FE99", x"FE9E", x"FEA5", x"FEAD", x"FEAB", x"FEBA", x"FEB1", x"FEAF", x"FEA7", x"FE9E", x"FE91", x"FE89", x"FE86", x"FE83", x"FE93", x"FEA8", x"FEC4", x"FEE9", x"FF0B", x"FF2C", x"FF40", x"FF5E", x"FF70", x"FF8A", x"FF9A", x"FFAC", x"FFAE", x"FFAF", x"FFAB", x"FFAA", x"FF9B", x"FF98", x"FF84", x"FF69", x"FF51", x"FF34", x"FF22", x"FF13", x"FF18", x"FF1A", x"FF21", x"FF30", x"FF32", x"FF39", x"FF39", x"FF32", x"FF2C", x"FF17", x"FF10", x"FEFD", x"FEF6", x"FEEE", x"FEE0", x"FEDD", x"FECF", x"FEC7", x"FEBA", x"FEB2", x"FEAA", x"FE9E", x"FEA4", x"FEA5", x"FEB6", x"FEC7", x"FEE3", x"FEEA", x"FEFB", x"FF01", x"FF09", x"FF13", x"FF1A", x"FF26", x"FF1B", x"FF21", x"FF1E", x"FF21", x"FF1E", x"FF25", x"FF11", x"FF0A", x"FEFA", x"FEF5", x"FEED", x"FEF2", x"FF03", x"FF0A", x"FF20", x"FF31", x"FF40", x"FF50", x"FF5F", x"FF70", x"FF81", x"FF94", x"FFAD", x"FFC0", x"FFD5", x"FFE9", x"FFF4", x"0001", x"FFFE", x"FFF7", x"FFE7", x"FFD2", x"FFC2", x"FFAD", x"FFB2", x"FFAD", x"FFBD", x"FFC5", x"FFD5", x"FFD4", x"FFD8", x"FFE0", x"FFDC", x"FFE6", x"FFE3", x"FFE4", x"FFD5", x"FFD1", x"FFCC", x"FFC9", x"FFCE", x"FFC9", x"FFC4", x"FFB1", x"FFA9", x"FFA0", x"FFA1", x"FFAC", x"FFC3", x"FFCF", x"FFE6", x"FFED", x"FFFB", x"FFFB", x"0004", x"0005", x"0009", x"000B", x"0004", x"0004", x"FFFB", x"FFF9", x"FFF2", x"FFE8", x"FFD5", x"FFBE", x"FFA6", x"FF8D", x"FF6D", x"FF5C", x"FF50", x"FF4C", x"FF58", x"FF71", x"FF7E", x"FF95", x"FFAB", x"FFC1", x"FFE4", x"0001", x"0027", x"0038", x"004D", x"005D", x"006D", x"0077", x"0089", x"008A", x"0086", x"007B", x"006B", x"005D", x"004C", x"004C", x"0046", x"004B", x"004D", x"004C", x"004A", x"0046", x"0044", x"003E", x"0041", x"003C", x"003E", x"0042", x"0044", x"004C", x"0041", x"0046", x"002C", x"0025", x"0016", x"000A", x"0000", x"0000", x"0004", x"0011", x"002C", x"004E", x"0068", x"0084", x"009D", x"00AA", x"00C0", x"00D0", x"00E3", x"00E4", x"00F2", x"00F4", x"00F8", x"00FB", x"00FC", x"00F8", x"00E6", x"00DC", x"00C6", x"00BC", x"00B7", x"00BB", x"00BB", x"00C3", x"00C6", x"00C2", x"00C3", x"00BC", x"00BA", x"00B0", x"00B2", x"00A4", x"00AC", x"00AC", x"00B7", x"00BD", x"00C6", x"00C9", x"00C3", x"00C3", x"00BF", x"00BD", x"00BA", x"00C3", x"00C6", x"00D2", x"00DE", x"00EA", x"00EB", x"00EF", x"00EE", x"00EF", x"00EC", x"00FC", x"00F6", x"00F8", x"00F7", x"00FA", x"0102", x"010B", x"0116", x"0113", x"010F", x"0109", x"0100", x"00F9", x"00FF", x"00F8", x"0105", x"00FD", x"0104", x"00FC", x"00F8", x"00F2", x"00ED", x"00EE", x"00EE", x"00F1", x"00F9", x"00FE", x"010A", x"010C", x"0117", x"010F", x"010E", x"0106", x"00FC", x"00F1", x"00E5", x"00E4", x"00DE", x"00E7", x"00F4", x"00FF", x"0100", x"0102", x"00F6", x"00F2", x"00EA", x"00EB", x"00E8", x"00E3", x"00E6", x"00E1", x"00E9", x"00ED", x"00F0", x"00F2", x"00EB", x"00ED", x"00EA", x"00EE", x"0102", x"0112", x"0132", x"0146", x"0158", x"0163", x"016A", x"0165", x"0169", x"0161", x"0160", x"015F", x"015B", x"0163", x"0156", x"0155", x"014C", x"013B", x"012C", x"0118", x"0105", x"00E8", x"00DC", x"00CC", x"00C9", x"00D5", x"00E8", x"00F0", x"0100", x"0105", x"010F", x"0118", x"0128", x"0134", x"013E", x"0145", x"014B", x"0153", x"0153", x"015F", x"0153", x"014B", x"0137", x"011F", x"0109", x"00FB", x"00F0", x"00F1", x"00EC", x"00F2", x"00E6", x"00E1", x"00E2", x"00D4", x"00DD", x"00DA", x"00DF", x"00DF", x"00EC", x"00F5", x"00FF", x"0107", x"010F", x"0109", x"010B", x"0106", x"00FF", x"0100", x"0104", x"0116", x"012C", x"0150", x"0170", x"018D", x"019E", x"01B4", x"01B9", x"01C8", x"01D1", x"01D0", x"01CF", x"01C6", x"01BE", x"01B3", x"01B0", x"01A9", x"019D", x"018B", x"017B", x"0167", x"0154", x"0153", x"014F", x"0155", x"015C", x"0162", x"0161", x"0162", x"0158", x"0149", x"013D", x"012D", x"0123", x"0119", x"0113", x"010D", x"0104", x"00FE", x"00F9", x"00EE", x"00E9", x"00DE", x"00D1", x"00C8", x"00C3", x"00C2", x"00CC", x"00D7", x"00E5", x"00F0", x"00F6", x"00FA", x"00F5", x"00F4", x"00F4", x"00F1", x"00F4", x"00F0", x"00F3", x"00EC", x"00EC", x"00E9", x"00E0", x"00E0", x"00D1", x"00CC", x"00C1", x"00C4", x"00C5", x"00D2", x"00DD", x"00F4", x"00F8", x"010D", x"010C", x"011A", x"011E", x"012C", x"0141", x"014F", x"016F", x"017C", x"0190", x"0195", x"0190", x"018B", x"0179", x"0169", x"0153", x"013F", x"0132", x"0122", x"0128", x"012A", x"0134", x"0134", x"0133", x"012B", x"011E", x"011C", x"0113", x"010B", x"0106", x"0101", x"00FA", x"00FE", x"0100", x"00FB", x"00F0", x"00E4", x"00D7", x"00D3", x"00DA", x"00E5", x"00F6", x"0109", x"0118", x"012C", x"0129", x"0137", x"0129", x"012E", x"0127", x"0126", x"0123", x"011C", x"011A", x"010F", x"010D", x"0101", x"00F2", x"00DF", x"00C4", x"00A8", x"0089", x"0076", x"0065", x"005A", x"0066", x"006F", x"0080", x"008F", x"00A1", x"00AA", x"00BC", x"00D1", x"00E1", x"00EE", x"00FE", x"010A", x"0110", x"0119", x"0122", x"0114", x"010C", x"00ED", x"00D5", x"00B1", x"00A0", x"0089", x"0082", x"0078", x"007B", x"0073", x"0074", x"0069", x"0062", x"0055", x"0051", x"004B", x"004D", x"0057", x"005C", x"0067", x"006D", x"006E", x"0067", x"0063", x"0054", x"0044", x"0032", x"0025", x"001E", x"0025", x"003F", x"0057", x"0077", x"008B", x"009A", x"00A0", x"00A1", x"00A9", x"00A6", x"00A6", x"00A7", x"00A3", x"00A4", x"00A0", x"009E", x"0090", x"0089", x"007B", x"0070", x"0067", x"0058", x"0058", x"0053", x"0060", x"0065", x"0071", x"006F", x"006C", x"0061", x"0055", x"004A", x"0044", x"0041", x"0045", x"0047", x"004F", x"0051", x"0059", x"0052", x"0056", x"004E", x"0047", x"0041", x"003E", x"0039", x"0040", x"004B", x"0055", x"0060", x"0064", x"0064", x"005B", x"0059", x"0054", x"004C", x"0044", x"0042", x"003A", x"003B", x"003B", x"003B", x"0035", x"0028", x"001E", x"0005", x"FFFC", x"FFE6", x"FFE1", x"FFD5", x"FFD0", x"FFCF", x"FFCC", x"FFCA", x"FFC9", x"FFC8", x"FFC6", x"FFCB", x"FFC6", x"FFD2", x"FFD6", x"FFE3", x"FFED", x"FFF9", x"FFF5", x"FFF5", x"FFE8", x"FFD6", x"FFBF", x"FFAD", x"FF98", x"FF91", x"FF90", x"FF9C", x"FFA7", x"FFAF", x"FFB5", x"FFB9", x"FFB1", x"FFBD", x"FFB4", x"FFB7", x"FFAE", x"FFB1", x"FFB0", x"FFB9", x"FFC4", x"FFC9", x"FFCE", x"FFCC", x"FFC8", x"FFC7", x"FFC3", x"FFCB", x"FFCE", x"FFDA", x"FFE5", x"FFE9", x"FFEE", x"FFE6", x"FFDF", x"FFD9", x"FFD0", x"FFCD", x"FFC7", x"FFC7", x"FFC1", x"FFBF", x"FFC1", x"FFB8", x"FFB1", x"FFA0", x"FF99", x"FF7C", x"FF70", x"FF55", x"FF43", x"FF39", x"FF3E", x"FF4E", x"FF61", x"FF71", x"FF83", x"FF83", x"FF8E", x"FF92", x"FF9F", x"FFA2", x"FFAF", x"FFB4", x"FFB7", x"FFBC", x"FFB8", x"FFAF", x"FF9E", x"FF89", x"FF71", x"FF59", x"FF42", x"FF31", x"FF23", x"FF1D", x"FF1B", x"FF1B", x"FF18", x"FF16", x"FF0A", x"FF0B", x"FEFD", x"FEFE", x"FEF7", x"FEFB", x"FEFF", x"FF06", x"FF16", x"FF14", x"FF19", x"FF14", x"FF13", x"FF09", x"FF08", x"FF07", x"FF0C", x"FF1D", x"FF3A", x"FF59", x"FF7D", x"FF9A", x"FFB2", x"FFBC", x"FFC4", x"FFC9", x"FFC6", x"FFC3", x"FFC2", x"FFB9", x"FFB6", x"FFAF", x"FFA6", x"FF9C", x"FF8E", x"FF7A", x"FF68", x"FF51", x"FF41", x"FF32", x"FF28", x"FF26", x"FF21", x"FF1E", x"FF19", x"FF09", x"FEFC", x"FEE3", x"FECC", x"FEB3", x"FE9A", x"FE8C", x"FE7D", x"FE7F", x"FE7D", x"FE7B", x"FE7A", x"FE7C", x"FE78", x"FE6D", x"FE6C", x"FE5C", x"FE5F", x"FE5E", x"FE73", x"FE7D", x"FE91", x"FE9D", x"FE9A", x"FE9C", x"FE98", x"FE98", x"FE95", x"FE96", x"FE98", x"FE91", x"FE9C", x"FE9D", x"FEAB", x"FEA6", x"FEB5", x"FEA6", x"FEA6", x"FE9D", x"FE98", x"FE95", x"FE98", x"FEA3", x"FEAC", x"FEBF", x"FECC", x"FED7", x"FEDF", x"FEE4", x"FEE9", x"FEEC", x"FEF5", x"FF04", x"FF0D", x"FF1E", x"FF2A", x"FF2F", x"FF36", x"FF2F", x"FF26", x"FF15", x"FF04", x"FEF2", x"FEE0", x"FEDF", x"FEDD", x"FEE3", x"FEEB", x"FEEE", x"FEE2", x"FEDF", x"FED5", x"FED0", x"FEC6", x"FEC8", x"FEBC", x"FEB8", x"FEB9", x"FEBC", x"FEBC", x"FEC4", x"FEBF", x"FEBE", x"FEB6", x"FEBD", x"FEBB", x"FEC1", x"FECC", x"FED0", x"FEDC", x"FEDF", x"FEEB", x"FEE6", x"FEEA", x"FEE3", x"FEDC", x"FED5", x"FEC8", x"FEC0", x"FEB1", x"FEA8", x"FE9A", x"FE91", x"FE7F", x"FE74", x"FE5B", x"FE4C", x"FE37", x"FE24", x"FE1B", x"FE1B", x"FE22", x"FE36", x"FE4A", x"FE60", x"FE6C", x"FE83", x"FE92", x"FEA6", x"FEBA", x"FECF", x"FEDB", x"FEE9", x"FEFA", x"FF01", x"FF03", x"FF02", x"FEF9", x"FEE9", x"FEDD", x"FED0", x"FEC2", x"FEB9", x"FEB1", x"FEB1", x"FEA9", x"FEAB", x"FEA5", x"FE9D", x"FE95", x"FE8B", x"FE84", x"FE7F", x"FE7B", x"FE79", x"FE7C", x"FE7E", x"FE82", x"FE82", x"FE78", x"FE6D", x"FE5C", x"FE51", x"FE46", x"FE40", x"FE4C", x"FE5A", x"FE77", x"FE9B", x"FEBB", x"FED1", x"FEDB", x"FEEE", x"FEED", x"FEFE", x"FEFC", x"FF02", x"FEF9", x"FEF5", x"FEF2", x"FEE3", x"FEDF", x"FED7", x"FEC9", x"FEBD", x"FEB3", x"FEB0", x"FEAB", x"FEAD", x"FEB8", x"FEBE", x"FECE", x"FED9", x"FEDE", x"FEDD", x"FED9", x"FECE", x"FEC8", x"FEBC", x"FEB9", x"FEB8", x"FEB5", x"FEBD", x"FEBF", x"FEC6", x"FECC", x"FED0", x"FED5", x"FED6", x"FED6", x"FED9", x"FEE4", x"FEF2", x"FF05", x"FF15", x"FF26", x"FF24", x"FF29", x"FF28", x"FF27", x"FF2A", x"FF2B", x"FF30", x"FF27", x"FF34", x"FF35", x"FF39", x"FF3E", x"FF3D", x"FF39", x"FF2E", x"FF2B", x"FF1A", x"FF12", x"FF01", x"FF02", x"FEF5", x"FF02", x"FF00", x"FF08", x"FF07", x"FF07", x"FF02", x"FF01", x"FEFD", x"FEFE", x"FF05", x"FF07", x"FF18", x"FF1A", x"FF23", x"FF1B", x"FF11", x"FF03", x"FEF2", x"FEDE", x"FED3", x"FECB", x"FEC4", x"FECF", x"FED6", x"FEDD", x"FEDF", x"FEDE", x"FEE2", x"FEDF", x"FEE8", x"FEEB", x"FEE9", x"FEF4", x"FEFB", x"FF0D", x"FF22", x"FF35", x"FF4D", x"FF53", x"FF64", x"FF69", x"FF76", x"FF81", x"FF8B", x"FF96", x"FF9B", x"FFA3", x"FFA4", x"FFA4", x"FFA4", x"FFA0", x"FF9D", x"FF95", x"FF92", x"FF7F", x"FF7A", x"FF69", x"FF5D", x"FF51", x"FF42", x"FF32", x"FF1F", x"FF0E", x"FEF6", x"FEE3", x"FED3", x"FED2", x"FED2", x"FEE3", x"FEF3", x"FEFB", x"FF09", x"FF11", x"FF26", x"FF37", x"FF59", x"FF6D", x"FF85", x"FF94", x"FFA3", x"FFAA", x"FFAE", x"FFAE", x"FF9E", x"FF8F", x"FF76", x"FF66", x"FF4A", x"FF3E", x"FF2B", x"FF24", x"FF1E", x"FF20", x"FF21", x"FF2B", x"FF36", x"FF41", x"FF53", x"FF5C", x"FF6D", x"FF73", x"FF86", x"FF8D", x"FF99", x"FFA4", x"FFA6", x"FFAC", x"FFAB", x"FFB1", x"FFB0", x"FFB5", x"FFC1", x"FFCF", x"FFE9", x"0004", x"0022", x"002E", x"003F", x"0047", x"004E", x"0057", x"005E", x"005E", x"005C", x"005E", x"0060", x"005D", x"0060", x"005D", x"004E", x"0044", x"0036", x"002C", x"0022", x"001F", x"001D", x"0017", x"001E", x"001D", x"001D", x"0019", x"0012", x"0002", x"FFF9", x"FFE7", x"FFDD", x"FFCE", x"FFC8", x"FFC5", x"FFBF", x"FFBD", x"FFC0", x"FFB5", x"FFBA", x"FFB1", x"FFB7", x"FFB0", x"FFC4", x"FFCA", x"FFE4", x"FFED", x"FFFE", x"FFF9", x"FFFD", x"FFF4", x"FFF6", x"FFF8", x"FFFC", x"0003", x"0006", x"000D", x"0019", x"001B", x"0029", x"0027", x"0027", x"0023", x"001E", x"0019", x"001A", x"001B", x"0022", x"0029", x"0039", x"0047", x"0056", x"0065", x"0074", x"007E", x"008B", x"009A", x"00A4", x"00B0", x"00BB", x"00C3", x"00CF", x"00D7", x"00DF", x"00DC", x"00DE", x"00CE", x"00C7", x"00B9", x"00B2", x"00A7", x"00A3", x"009E", x"0092", x"0085", x"007C", x"006B", x"006A", x"0061", x"0067", x"005E", x"0067", x"006B", x"007C", x"008D", x"00A8", x"00BA", x"00BF", x"00D1", x"00CC", x"00D6", x"00D9", x"00E4", x"00E1", x"00E3", x"00E7", x"00DE", x"00E0", x"00DE", x"00DA", x"00D4", x"00CD", x"00C5", x"00B7", x"00B0", x"00A5", x"00A0", x"009D", x"0098", x"0095", x"008B", x"0086", x"0076", x"006C", x"0068", x"0063", x"006A", x"007B", x"008B", x"009A", x"00A6", x"00B4", x"00BC", x"00D1", x"00E0", x"00F7", x"00FC", x"0114", x"0119", x"011F", x"012B", x"0122", x"011D", x"00FF", x"00F7", x"00DB", x"00D3", x"00CB", x"00BE", x"00B2", x"00A7", x"009F", x"009A", x"0099", x"009B", x"009F", x"00A5", x"00AF", x"00B9", x"00C4", x"00C9", x"00D3", x"00D3", x"00D8", x"00D4", x"00CD", x"00C5", x"00B6", x"00AB", x"00A5", x"00A4", x"00AD", x"00B7", x"00D2", x"00E2", x"00FC", x"010A", x"011D", x"0126", x"0131", x"0142", x"0141", x"0143", x"0146", x"013D", x"013D", x"0142", x"013B", x"0136", x"012A", x"0124", x"0115", x"0117", x"0115", x"0118", x"0115", x"0118", x"011C", x"011B", x"0122", x"0122", x"0122", x"0120", x"011C", x"0116", x"010A", x"0106", x"00FC", x"00FD", x"0102", x"0106", x"0110", x"0114", x"0119", x"011D", x"0122", x"012F", x"0137", x"014D", x"015E", x"0168", x"016E", x"016D", x"0163", x"015C", x"015C", x"0159", x"0153", x"014C", x"014B", x"0140", x"0148", x"0148", x"0146", x"0133", x"0127", x"0110", x"0103", x"00F6", x"00F1", x"00EA", x"00E7", x"00EB", x"00F0", x"00F7", x"0105", x"010D", x"0115", x"0119", x"011E", x"011C", x"011E", x"011B", x"011B", x"0119", x"0116", x"010A", x"0103", x"00F5", x"00E7", x"00DB", x"00D8", x"00CC", x"00CF", x"00D7", x"00DE", x"00E6", x"00E9", x"00F0", x"00EC", x"00F0", x"00FC", x"00F8", x"00FD", x"0105", x"010E", x"011F", x"013B", x"0158", x"0166", x"0174", x"0180", x"0181", x"018C", x"0196", x"019D", x"019D", x"019C", x"0196", x"018F", x"0189", x"018E", x"0186", x"0189", x"0182", x"0173", x"0168", x"0156", x"0148", x"0136", x"0127", x"0120", x"010B", x"0108", x"00FA", x"00EA", x"00DE", x"00D0", x"00C3", x"00BC", x"00C6", x"00C0", x"00C9", x"00C5", x"00CE", x"00D1", x"00E3", x"00F7", x"0104", x"011A", x"0125", x"013A", x"0142", x"0159", x"015C", x"014F", x"0143", x"0128", x"010C", x"00F7", x"00DC", x"00D1", x"00B5", x"00B6", x"00A3", x"00AC", x"00AB", x"00BD", x"00C6", x"00D8", x"00E8", x"00ED", x"00FC", x"00FA", x"0100", x"0100", x"0105", x"0107", x"010A", x"0109", x"010E", x"0106", x"010C", x"010C", x"0112", x"012A", x"013B", x"0155", x"0164", x"0178", x"017F", x"0186", x"018F", x"018A", x"018E", x"0182", x"0185", x"0175", x"0170", x"0168", x"0155", x"0144", x"012A", x"0112", x"00F7", x"00E8", x"00D8", x"00CD", x"00BE", x"00B4", x"00A0", x"0099", x"0092", x"008A", x"008A", x"007F", x"007A", x"006B", x"0060", x"0056", x"004A", x"0046", x"003F", x"003D", x"0035", x"003B", x"002D", x"002F", x"002C", x"0020", x"0029", x"0025", x"0030", x"0032", x"0036", x"003B", x"003A", x"0041", x"004E", x"0058", x"0061", x"0070", x"0070", x"0073", x"007C", x"007F", x"007B", x"0079", x"006F", x"0061", x"0060", x"005C", x"0062", x"0063", x"0065", x"0069", x"006A", x"0073", x"0084", x"0088", x"009A", x"009C", x"00A1", x"009C", x"00A1", x"0094", x"0098", x"0092", x"0097", x"0095", x"0096", x"0095", x"008D", x"0086", x"007C", x"0074", x"0069", x"0069", x"0058", x"0053", x"0045", x"0034", x"002B", x"001D", x"001A", x"0013", x"0011", x"0018", x"0013", x"0026", x"002E", x"0046", x"0051", x"0060", x"0062", x"005D", x"0063", x"0062", x"0063", x"0067", x"0062", x"005B", x"004A", x"0047", x"0039", x"0034", x"0032", x"0026", x"001C", x"000E", x"0001", x"FFF3", x"FFE6", x"FFD9", x"FFD5", x"FFC4", x"FFC8", x"FFB9", x"FFB4", x"FFAE", x"FFA3", x"FF9E", x"FF99", x"FFA5", x"FFA5", x"FFB7", x"FFBE", x"FFC7", x"FFD2", x"FFE9", x"FFFA", x"0015", x"0025", x"003D", x"0042", x"0052", x"0059", x"0057", x"0050", x"0042", x"0025", x"0011", x"FFF8", x"FFE8", x"FFD0", x"FFC0", x"FFA6", x"FF8E", x"FF77", x"FF71", x"FF63", x"FF64", x"FF65", x"FF66", x"FF6A", x"FF6A", x"FF69", x"FF64", x"FF60", x"FF5C", x"FF59", x"FF53", x"FF54", x"FF47", x"FF4D", x"FF42", x"FF44", x"FF44", x"FF4C", x"FF58", x"FF67", x"FF7C", x"FF87", x"FF8E", x"FF91", x"FF95", x"FF94", x"FF96", x"FF99", x"FF94", x"FF93", x"FF99", x"FF99", x"FF9D", x"FF9D", x"FF95", x"FF8A", x"FF7B", x"FF7F", x"FF74", x"FF74", x"FF74", x"FF69", x"FF65", x"FF64", x"FF6B", x"FF72", x"FF82", x"FF87", x"FF85", x"FF7D", x"FF73", x"FF5D", x"FF53", x"FF44", x"FF40", x"FF3B", x"FF3F", x"FF45", x"FF46", x"FF4C", x"FF52", x"FF54", x"FF5E", x"FF6A", x"FF6E", x"FF7B", x"FF78", x"FF77", x"FF69", x"FF68", x"FF6A", x"FF6A", x"FF77", x"FF76", x"FF7A", x"FF71", x"FF7D", x"FF71", x"FF75", x"FF66", x"FF58", x"FF3C", x"FF2E", x"FF22", x"FF16", x"FF13", x"FF0E", x"FF04", x"FF01", x"FF00", x"FF08", x"FF0B", x"FF19", x"FF1F", x"FF22", x"FF24", x"FF25", x"FF1A", x"FF14", x"FF07", x"FF00", x"FEF7", x"FEF5", x"FEF2", x"FEE6", x"FEE2", x"FEDF", x"FECE", x"FED8", x"FECE", x"FED0", x"FECD", x"FEC5", x"FEBD", x"FEAE", x"FEAE", x"FEA9", x"FEAE", x"FEB3", x"FEBC", x"FEC7", x"FED2", x"FEED", x"FEF9", x"FF14", x"FF27", x"FF34", x"FF43", x"FF4E", x"FF5B", x"FF63", x"FF6A", x"FF6D", x"FF64", x"FF5F", x"FF51", x"FF4B", x"FF3D", x"FF3D", x"FF27", x"FF1F", x"FF07", x"FEF3", x"FED9", x"FEC6", x"FEB2", x"FEA3", x"FE98", x"FE93", x"FE87", x"FE82", x"FE76", x"FE6A", x"FE5A", x"FE54", x"FE4A", x"FE48", x"FE4C", x"FE4F", x"FE4D", x"FE59", x"FE65", x"FE79", x"FE98", x"FEB3", x"FED0", x"FEE0", x"FEFC", x"FF04", x"FF10", x"FF06", x"FEFE", x"FED9", x"FEC4", x"FEA7", x"FE95", x"FE87", x"FE7D", x"FE77", x"FE67", x"FE6D", x"FE6E", x"FE79", x"FE86", x"FE9C", x"FEA9", x"FEBB", x"FECC", x"FED1", x"FEDD", x"FEDE", x"FEE2", x"FEE6", x"FEED", x"FEF5", x"FEF4", x"FEF7", x"FEF3", x"FEF2", x"FEF9", x"FF03", x"FF17", x"FF21", x"FF39", x"FF39", x"FF43", x"FF40", x"FF45", x"FF47", x"FF4A", x"FF4B", x"FF48", x"FF3F", x"FF40", x"FF38", x"FF33", x"FF2F", x"FF26", x"FF18", x"FF13", x"FF05", x"FF09", x"FEFB", x"FEFF", x"FEED", x"FEDE", x"FED5", x"FEC3", x"FEC1", x"FEBC", x"FEBB", x"FEB4", x"FEAF", x"FEA1", x"FE92", x"FE83", x"FE79", x"FE74", x"FE74", x"FE7B", x"FE83", x"FE86", x"FE8F", x"FE8E", x"FE8D", x"FE90", x"FE96", x"FE9C", x"FEA8", x"FEB0", x"FEB3", x"FEB5", x"FEC0", x"FEC9", x"FEDD", x"FEEA", x"FEFD", x"FEF8", x"FF04", x"FEFB", x"FF00", x"FEFC", x"FEFB", x"FEF4", x"FEE5", x"FEE6", x"FED9", x"FEE3", x"FEDC", x"FEE9", x"FEE7", x"FEF0", x"FEFB", x"FF03", x"FF16", x"FF22", x"FF33", x"FF3C", x"FF47", x"FF44", x"FF44", x"FF3A", x"FF31", x"FF2A", x"FF22", x"FF22", x"FF1D", x"FF18", x"FF19", x"FF0E", x"FF11", x"FF0A", x"FF0B", x"FF04", x"FEFB", x"FEF3", x"FEDA", x"FECF", x"FEBF", x"FEBC", x"FEBD", x"FEC8", x"FED3", x"FEE0", x"FEF6", x"FF11", x"FF28", x"FF49", x"FF60", x"FF74", x"FF80", x"FF8E", x"FF98", x"FF9D", x"FFA3", x"FF9D", x"FF93", x"FF86", x"FF77", x"FF6A", x"FF65", x"FF5D", x"FF5E", x"FF5E", x"FF59", x"FF57", x"FF43", x"FF3E", x"FF2F", x"FF29", x"FF2B", x"FF2A", x"FF2C", x"FF33", x"FF32", x"FF34", x"FF32", x"FF39", x"FF37", x"FF40", x"FF44", x"FF45", x"FF45", x"FF4D", x"FF58", x"FF69", x"FF83", x"FF9E", x"FFAB", x"FFBE", x"FFC3", x"FFCB", x"FFCB", x"FFC8", x"FFBD", x"FFA6", x"FF91", x"FF77", x"FF64", x"FF52", x"FF47", x"FF3A", x"FF2F", x"FF25", x"FF24", x"FF1E", x"FF2D", x"FF2F", x"FF3F", x"FF47", x"FF53", x"FF55", x"FF55", x"FF57", x"FF50", x"FF50", x"FF51", x"FF52", x"FF53", x"FF52", x"FF53", x"FF4C", x"FF52", x"FF5F", x"FF66", x"FF80", x"FF89", x"FF95", x"FF99", x"FF9F", x"FFAA", x"FFB2", x"FFBF", x"FFCE", x"FFCE", x"FFDA", x"FFDF", x"FFE6", x"FFE8", x"FFED", x"FFE9", x"FFE1", x"FFDB", x"FFD7", x"FFCD", x"FFCC", x"FFC4", x"FFC4", x"FFBF", x"FFC4", x"FFC8", x"FFD2", x"FFDD", x"FFEC", x"FFF4", x"FFFC", x"FFF6", x"FFF2", x"FFE4", x"FFDF", x"FFD6", x"FFDB", x"FFDB", x"FFE3", x"FFE9", x"FFF4", x"FFF8", x"0002", x"0008", x"0012", x"0011", x"001F", x"0015", x"0014", x"0009", x"0008", x"0006", x"000D", x"0010", x"001B", x"0010", x"0019", x"000C", x"000D", x"000A", x"0007", x"0000", x"FFF1", x"FFEB", x"FFDF", x"FFDC", x"FFDE", x"FFE2", x"FFDE", x"FFE8", x"FFE7", x"FFEC", x"FFF5", x"FFFC", x"0003", x"000D", x"000C", x"000F", x"0008", x"0005", x"0001", x"FFFC", x"0000", x"0002", x"0006", x"000F", x"0016", x"0018", x"0019", x"001E", x"001B", x"0020", x"001E", x"001A", x"000F", x"000A", x"0005", x"000D", x"0017", x"002B", x"0033", x"0041", x"004F", x"005E", x"0071", x"008A", x"009D", x"00B0", x"00BA", x"00CC", x"00D2", x"00DD", x"00E1", x"00E1", x"00D7", x"00D3", x"00C4", x"00BD", x"00B3", x"00AE", x"00AC", x"00A7", x"00A8", x"009A", x"0095", x"0089", x"007C", x"0077", x"0072", x"006B", x"006D", x"0066", x"0060", x"0053", x"004A", x"003E", x"0037", x"002F", x"0031", x"0027", x"0026", x"0028", x"0031", x"0043", x"005E", x"007F", x"0093", x"00B0", x"00BE", x"00CD", x"00D4", x"00DB", x"00D2", x"00C4", x"00B2", x"009B", x"0086", x"0079", x"0070", x"0065", x"005E", x"005D", x"005A", x"0061", x"0067", x"0079", x"0084", x"0099", x"00A6", x"00B6", x"00C2", x"00CE", x"00D3", x"00DF", x"00E4", x"00ED", x"00F3", x"00FD", x"0101", x"0104", x"0111", x"0116", x"0127", x"0133", x"013B", x"013C", x"0139", x"0137", x"0133", x"013A", x"013F", x"0146", x"013D", x"013C", x"0133", x"0124", x"0123", x"0116", x"010B", x"00FE", x"00EE", x"00E4", x"00D4", x"00CA", x"00C1", x"00AF", x"00A7", x"009B", x"0095", x"0091", x"0095", x"0093", x"0096", x"0097", x"0092", x"008B", x"0084", x"0079", x"0074", x"006B", x"006E", x"006C", x"006D", x"0076", x"006E", x"0074", x"0073", x"007A", x"0084", x"0094", x"009D", x"00A6", x"00AF", x"00B9", x"00C4", x"00D7", x"00E6", x"00EF", x"00F6", x"00F2", x"00F9", x"00F3", x"00FB", x"00F9", x"00F4", x"00F1", x"00E7", x"00E1", x"00DC", x"00DD", x"00DD", x"00E0", x"00E5", x"00EF", x"00F4", x"0101", x"0108", x"010E", x"0116", x"0119", x"011A", x"0115", x"0118", x"010B", x"0108", x"0105", x"0102", x"0107", x"0112", x"0116", x"011C", x"011A", x"011E", x"0117", x"0115", x"0111", x"00FE", x"00E7", x"00D2", x"00B9", x"00A8", x"00A6", x"00A8", x"00AB", x"00B6", x"00C7", x"00D6", x"00F7", x"0112", x"0132", x"0149", x"015B", x"0170", x"0179", x"0182", x"0188", x"017C", x"0174", x"0166", x"0153", x"0149", x"013B", x"0138", x"012D", x"012C", x"0125", x"011E", x"0114", x"010B", x"00F9", x"00F3", x"00E7", x"00E7", x"00E3", x"00E7", x"00E0", x"00D7", x"00D1", x"00C6", x"00BF", x"00C0", x"00C4", x"00C1", x"00CB", x"00CF", x"00E0", x"00F2", x"0117", x"012C", x"0149", x"0155", x"0166", x"0163", x"0164", x"0160", x"014E", x"013A", x"0124", x"0103", x"00EB", x"00D0", x"00BE", x"00A5", x"0096", x"0085", x"0081", x"0076", x"007C", x"007D", x"007F", x"008B", x"008F", x"009A", x"00A1", x"00A8", x"00AA", x"00B2", x"00B5", x"00BA", x"00C1", x"00C4", x"00C9", x"00C5", x"00C7", x"00C9", x"00C9", x"00D8", x"00D8", x"00E0", x"00DC", x"00E1", x"00DF", x"00E8", x"00F7", x"00FC", x"010C", x"0110", x"011B", x"011A", x"0122", x"011E", x"011E", x"0110", x"010C", x"00F7", x"00F1", x"00DF", x"00DA", x"00CF", x"00CB", x"00CB", x"00C8", x"00CE", x"00CE", x"00D5", x"00D2", x"00D8", x"00D1", x"00CE", x"00CB", x"00C0", x"00BC", x"00B7", x"00B0", x"00B1", x"00B2", x"00B9", x"00B5", x"00BB", x"00C0", x"00C0", x"00CD", x"00D4", x"00E0", x"00DE", x"00E4", x"00E3", x"00E6", x"00EB", x"00FC", x"00F6", x"00F7", x"00EE", x"00E8", x"00DE", x"00D8", x"00D0", x"00BD", x"00B1", x"00A3", x"0099", x"0090", x"0095", x"0092", x"0095", x"009A", x"00A1", x"00A4", x"00A6", x"00A6", x"00A3", x"00A6", x"00A3", x"00A9", x"00A1", x"00A0", x"0098", x"0094", x"009B", x"0095", x"00A5", x"00A1", x"00A9", x"00A0", x"009C", x"0092", x"0086", x"0083", x"0077", x"0071", x"0058", x"0052", x"0036", x"0032", x"0031", x"0033", x"003A", x"0040", x"004D", x"005C", x"0077", x"0095", x"00AE", x"00C8", x"00D7", x"00E9", x"00E8", x"00F1", x"00EC", x"00E5", x"00DA", x"00CE", x"00B9", x"00AA", x"0096", x"0082", x"006E", x"0061", x"004B", x"003F", x"002F", x"0025", x"0014", x"000D", x"0004", x"0001", x"FFF9", x"FFFD", x"FFED", x"FFE6", x"FFD7", x"FFC6", x"FFBF", x"FFBA", x"FFBF", x"FFB5", x"FFB8", x"FFB6", x"FFBB", x"FFC4", x"FFE0", x"FFF3", x"000E", x"0023", x"0035", x"0041", x"004D", x"0057", x"0052", x"004D", x"0040", x"002D", x"0019", x"000A", x"FFFD", x"FFEB", x"FFE6", x"FFD9", x"FFD8", x"FFD5", x"FFDE", x"FFE1", x"FFF0", x"FFFC", x"000C", x"001E", x"002E", x"0040", x"0049", x"0056", x"005A", x"005C", x"0061", x"005E", x"0059", x"0051", x"004B", x"003F", x"003D", x"003B", x"0037", x"0032", x"0029", x"0025", x"0022", x"0024", x"0032", x"0030", x"0040", x"003D", x"0045", x"0043", x"004A", x"004A", x"0043", x"003C", x"002D", x"0018", x"0007", x"FFF2", x"FFE5", x"FFCF", x"FFCA", x"FFBE", x"FFB2", x"FFB2", x"FFA8", x"FFA5", x"FFA0", x"FF9A", x"FF95", x"FF95", x"FF88", x"FF8C", x"FF79", x"FF80", x"FF73", x"FF72", x"FF75", x"FF6B", x"FF6E", x"FF66", x"FF69", x"FF65", x"FF6D", x"FF78", x"FF7A", x"FF89", x"FF89", x"FF8A", x"FF8F", x"FF96", x"FFA2", x"FFA5", x"FFA9", x"FFA7", x"FFA1", x"FF9C", x"FF9D", x"FF97", x"FF90", x"FF86", x"FF80", x"FF72", x"FF70", x"FF71", x"FF6C", x"FF72", x"FF7C", x"FF82", x"FF8A", x"FF93", x"FF92", x"FF8F", x"FF89", x"FF85", x"FF7C", x"FF7A", x"FF72", x"FF67", x"FF5C", x"FF53", x"FF4C", x"FF45", x"FF41", x"FF3A", x"FF30", x"FF2A", x"FF1E", x"FF18", x"FF12", x"FF11", x"FF09", x"FEFF", x"FEF2", x"FEDE", x"FED7", x"FED4", x"FEDB", x"FEE3", x"FEF5", x"FF0A", x"FF20", x"FF41", x"FF63", x"FF7F", x"FF9D", x"FFAE", x"FFBF", x"FFC3", x"FFCB", x"FFCA", x"FFBF", x"FFBC", x"FFAB", x"FFA1", x"FF8F", x"FF84", x"FF71", x"FF5F", x"FF53", x"FF3E", x"FF39", x"FF2D", x"FF2B", x"FF22", x"FF25", x"FF20", x"FF1C", x"FF21", x"FF19", x"FF1B", x"FF0D", x"FF07", x"FEF7", x"FEEA", x"FEEC", x"FEE1", x"FEDF", x"FEDB", x"FED7", x"FED8", x"FEE4", x"FEF7", x"FF09", x"FF1B", x"FF2D", x"FF32", x"FF3E", x"FF41", x"FF4B", x"FF42", x"FF3F", x"FF2D", x"FF1C", x"FF03", x"FEF5", x"FEDF", x"FECC", x"FEBD", x"FEAB", x"FEA2", x"FE98", x"FE98", x"FE90", x"FE8C", x"FE8F", x"FE89", x"FE91", x"FE9F", x"FEA2", x"FEB9", x"FEBB", x"FECD", x"FECE", x"FED7", x"FED3", x"FECE", x"FEC2", x"FEBB", x"FEAD", x"FEAF", x"FEB2", x"FEB9", x"FEB8", x"FEC2", x"FEBC", x"FEC1", x"FECB", x"FED7", x"FEE9", x"FEF8", x"FF0C", x"FF11", x"FF20", x"FF2D", x"FF30", x"FF33", x"FF2B", x"FF1C", x"FF07", x"FEF9", x"FEEB", x"FED8", x"FED4", x"FECE", x"FECE", x"FED5", x"FED8", x"FEE1", x"FEE0", x"FEE4", x"FEE9", x"FEE8", x"FEF4", x"FEF5", x"FEF9", x"FEF9", x"FEF3", x"FEF2", x"FEE3", x"FEE5", x"FED8", x"FED3", x"FECA", x"FEC4", x"FEBE", x"FEC4", x"FEC9", x"FED1", x"FED3", x"FED7", x"FED5", x"FED4", x"FEDC", x"FEE2", x"FEE5", x"FEEE", x"FEE7", x"FEE6", x"FEE0", x"FEE0", x"FED9", x"FED3", x"FECF", x"FEBF", x"FEBE", x"FEAF", x"FEB3", x"FEA5", x"FEAA", x"FEA9", x"FEA5", x"FEAD", x"FEAB", x"FEA7", x"FEA2", x"FE94", x"FE8E", x"FE81", x"FE83", x"FE82", x"FE87", x"FE91", x"FE9E", x"FEA6", x"FEB3", x"FEBF", x"FEC0", x"FEC2", x"FEBF", x"FEB3", x"FEB3", x"FEB3", x"FEB7", x"FEB0", x"FEAF", x"FEA9", x"FE9A", x"FE9A", x"FE9A", x"FEA1", x"FEA4", x"FEB5", x"FEC4", x"FED7", x"FEF9", x"FF14", x"FF35", x"FF47", x"FF61", x"FF65", x"FF70", x"FF75", x"FF76", x"FF77", x"FF74", x"FF75", x"FF68", x"FF66", x"FF59", x"FF45", x"FF3A", x"FF25", x"FF14", x"FF01", x"FEFF", x"FEF3", x"FEEF", x"FEEF", x"FEE1", x"FEDC", x"FED0", x"FEC8", x"FEB8", x"FEAB", x"FE9D", x"FE8C", x"FE83", x"FE87", x"FE81", x"FE88", x"FE82", x"FE88", x"FE80", x"FE94", x"FE9F", x"FEB6", x"FEC9", x"FEDD", x"FEF1", x"FEFF", x"FF15", x"FF22", x"FF25", x"FF2D", x"FF26", x"FF1C", x"FF15", x"FF08", x"FEFD", x"FEF3", x"FEEC", x"FEE4", x"FEE1", x"FEE9", x"FEE5", x"FEEB", x"FEEF", x"FEF4", x"FEFB", x"FF0F", x"FF27", x"FF3F", x"FF5F", x"FF72", x"FF8A", x"FF95", x"FFA7", x"FFAC", x"FFAB", x"FFA9", x"FF9D", x"FF89", x"FF88", x"FF7B", x"FF7E", x"FF7A", x"FF7A", x"FF72", x"FF69", x"FF69", x"FF63", x"FF69", x"FF6B", x"FF78", x"FF76", x"FF80", x"FF87", x"FF89", x"FF86", x"FF88", x"FF76", x"FF6F", x"FF5F", x"FF56", x"FF47", x"FF43", x"FF3E", x"FF3D", x"FF3D", x"FF43", x"FF3D", x"FF3E", x"FF35", x"FF2D", x"FF21", x"FF23", x"FF1E", x"FF26", x"FF25", x"FF2C", x"FF20", x"FF23", x"FF1C", x"FF1A", x"FF12", x"FF13", x"FF0D", x"FF14", x"FF1D", x"FF35", x"FF42", x"FF59", x"FF65", x"FF70", x"FF75", x"FF83", x"FF84", x"FF95", x"FF93", x"FFA1", x"FF9E", x"FFA6", x"FFAD", x"FFAE", x"FFB4", x"FFB0", x"FFA8", x"FF9F", x"FF98", x"FF92", x"FF8E", x"FF92", x"FF92", x"FF99", x"FFA0", x"FFA8", x"FFA7", x"FFAA", x"FFA3", x"FF9E", x"FF97", x"FF9D", x"FF9E", x"FFA8", x"FFB2", x"FFBA", x"FFBD", x"FFCA", x"FFC9", x"FFCD", x"FFC7", x"FFBF", x"FFB6", x"FFAA", x"FFAE", x"FFA8", x"FFAA", x"FFA9", x"FFA2", x"FF99", x"FF9A", x"FF99", x"FFA1", x"FFB0", x"FFBF", x"FFD9", x"FFF0", x"0017", x"003B", x"0059", x"007B", x"008E", x"00A0", x"00A7", x"00B5", x"00AA", x"00B1", x"00A8", x"00A1", x"009E", x"0090", x"008B", x"0074", x"0062", x"004C", x"002F", x"0024", x"0013", x"0011", x"000B", x"000F", x"000C", x"000C", x"000F", x"0011", x"0014", x"0013", x"0017", x"0008", x"0011", x"000B", x"0019", x"0027", x"0033", x"0041", x"0044", x"0051", x"0059", x"0066", x"0071", x"0081", x"0086", x"0098", x"009F", x"00AF", x"00AE", x"00B2", x"00A3", x"0090", x"0084", x"0068", x"0055", x"0044", x"002F", x"0023", x"0019", x"0017", x"000F", x"000D", x"000B", x"0006", x"0005", x"0010", x"0019", x"002D", x"0043", x"0057", x"0064", x"0072", x"007E", x"0080", x"007E", x"0075", x"006A", x"0058", x"0059", x"0051", x"0059", x"005C", x"0068", x"005F", x"0068", x"0069", x"0075", x"0083", x"009B", x"00A8", x"00BC", x"00D3", x"00E7", x"00F6", x"00FF", x"0108", x"00FA", x"00F0", x"00E6", x"00D5", x"00CC", x"00C4", x"00BB", x"00B7", x"00B3", x"00BA", x"00B1", x"00B5", x"00B2", x"00B0", x"00AF", x"00B6", x"00B9", x"00C0", x"00C8", x"00CF", x"00D5", x"00D8", x"00DB", x"00D7", x"00D5", x"00D1", x"00C8", x"00CA", x"00CD", x"00D9", x"00E6", x"00F7", x"00FF", x"0103", x"0105", x"010A", x"0103", x"010F", x"0108", x"0108", x"0101", x"0108", x"0100", x"010C", x"010B", x"010D", x"0100", x"00FD", x"00F2", x"00EB", x"00E8", x"00E7", x"00E0", x"00E5", x"00E5", x"00EB", x"00E7", x"00E4", x"00DB", x"00CB", x"00C2", x"00C6", x"00BF", x"00D3", x"00DC", x"00EE", x"00F2", x"0102", x"0100", x"00FE", x"00FB", x"00EB", x"00DF", x"00D2", x"00CC", x"00CB", x"00CF", x"00CF", x"00D4", x"00C8", x"00CD", x"00C5", x"00C8", x"00CC", x"00D8", x"00E6", x"0101", x"0127", x"013F", x"0165", x"0178", x"0189", x"018B", x"0195", x"0191", x"0190", x"0188", x"0183", x"0172", x"016E", x"015D", x"0154", x"013E", x"0129", x"0112", x"00F9", x"00E8", x"00DF", x"00D2", x"00D7", x"00D1", x"00D6", x"00D5", x"00D3", x"00CF", x"00C7", x"00C3", x"00B1", x"00AD", x"009C", x"009D", x"009C", x"00A4", x"00AE", x"00AD", x"00B2", x"00B3", x"00B0", x"00BF", x"00C6", x"00D1", x"00DB", x"00EF", x"00FE", x"0113", x"0120", x"0135", x"0123", x"012A", x"0118", x"0112", x"0100", x"00FA", x"00E9", x"00E2", x"00DD", x"00E0", x"00E2", x"00E4", x"00ED", x"00E8", x"00EF", x"00F8", x"0108", x"0116", x"012F", x"0143", x"0159", x"016F", x"017D", x"0185", x"0181", x"0173", x"0160", x"0149", x"013D", x"0132", x"0131", x"0133", x"0137", x"0134", x"0135", x"0130", x"012F", x"012D", x"0133", x"012F", x"0135", x"013D", x"0140", x"014C", x"014D", x"014D", x"0138", x"012F", x"0119", x"0104", x"00F7", x"00E6", x"00DE", x"00CF", x"00D6", x"00CE", x"00D3", x"00D1", x"00CC", x"00C9", x"00BF", x"00BF", x"00C0", x"00C2", x"00CC", x"00CD", x"00D6", x"00D3", x"00D3", x"00C8", x"00BD", x"00B3", x"00A5", x"00A3", x"00A3", x"00A6", x"00B5", x"00BF", x"00CC", x"00D0", x"00D8", x"00D6", x"00D8", x"00DE", x"00DD", x"00E2", x"00E9", x"00F1", x"00F7", x"0103", x"0107", x"0108", x"0101", x"00FD", x"00F5", x"00EE", x"00E8", x"00E6", x"00D5", x"00DA", x"00D2", x"00D1", x"00CA", x"00C8", x"00B3", x"00A7", x"0094", x"008E", x"0082", x"0083", x"0087", x"0087", x"008D", x"0092", x"008D", x"008E", x"0083", x"0075", x"0066", x"0053", x"004F", x"0041", x"0048", x"0048", x"004C", x"004C", x"0052", x"0050", x"0056", x"0060", x"0067", x"0078", x"008C", x"00AC", x"00C7", x"00EC", x"0103", x"0119", x"0117", x"0128", x"011C", x"011E", x"0117", x"0111", x"0107", x"0105", x"0100", x"00F8", x"00E7", x"00D7", x"00C0", x"00A9", x"0099", x"0088", x"0082", x"007E", x"0080", x"0087", x"0090", x"0094", x"0092", x"008D", x"007A", x"006A", x"0053", x"0046", x"003D", x"003D", x"004B", x"004C", x"0054", x"005A", x"0055", x"005A", x"005D", x"0066", x"006C", x"0077", x"0086", x"0094", x"00A4", x"00B6", x"00B9", x"00B2", x"00A0", x"0091", x"006F", x"005E", x"0044", x"002C", x"001B", x"0009", x"0000", x"FFF1", x"FFF0", x"FFE3", x"FFE4", x"FFDA", x"FFE1", x"FFE1", x"FFEC", x"FFFF", x"0012", x"0028", x"003B", x"0047", x"004A", x"004C", x"003E", x"002D", x"0018", x"0003", x"FFFC", x"FFF2", x"FFFD", x"FFFA", x"FFFE", x"0002", x"0000", x"0007", x"0009", x"000A", x"000E", x"000D", x"001B", x"0023", x"0034", x"0046", x"0049", x"0048", x"0046", x"0035", x"0028", x"0018", x"0006", x"FFF9", x"FFED", x"FFEF", x"FFF0", x"FFF4", x"FFF8", x"FFFB", x"FFF1", x"FFF6", x"FFE8", x"FFEB", x"FFE9", x"FFF0", x"FFF3", x"FFFF", x"0000", x"0005", x"FFFA", x"FFF4", x"FFE5", x"FFCF", x"FFC4", x"FFB7", x"FFAF", x"FFBB", x"FFBF", x"FFCC", x"FFD5", x"FFDD", x"FFDA", x"FFE1", x"FFD8", x"FFE0", x"FFD6", x"FFDE", x"FFE0", x"FFE8", x"FFF1", x"FFF8", x"FFF8", x"FFED", x"FFEA", x"FFD6", x"FFCB", x"FFB9", x"FFB2", x"FFA1", x"FFA3", x"FF9D", x"FF9E", x"FF96", x"FF96", x"FF86", x"FF81", x"FF75", x"FF70", x"FF6E", x"FF77", x"FF7C", x"FF8A", x"FF95", x"FFA2", x"FFA4", x"FFAF", x"FFA6", x"FF9E", x"FF91", x"FF80", x"FF74", x"FF69", x"FF6C", x"FF67", x"FF64", x"FF62", x"FF59", x"FF54", x"FF52", x"FF55", x"FF54", x"FF5A", x"FF6A", x"FF7C", x"FF99", x"FFBA", x"FFD7", x"FFEC", x"FFF8", x"0005", x"0000", x"FFFE", x"FFFC", x"FFEE", x"FFEB", x"FFDC", x"FFD5", x"FFC4", x"FFB6", x"FFA0", x"FF89", x"FF70", x"FF5F", x"FF47", x"FF3E", x"FF36", x"FF31", x"FF31", x"FF35", x"FF34", x"FF37", x"FF37", x"FF2B", x"FF1F", x"FF0F", x"FEFC", x"FEF9", x"FEF3", x"FF03", x"FF03", x"FF0E", x"FF12", x"FF15", x"FF14", x"FF18", x"FF1D", x"FF1C", x"FF29", x"FF31", x"FF41", x"FF56", x"FF66", x"FF70", x"FF6F", x"FF67", x"FF54", x"FF3F", x"FF28", x"FF18", x"FF07", x"FEFE", x"FEFD", x"FEFD", x"FF03", x"FF07", x"FF0E", x"FF0D", x"FF17", x"FF14", x"FF24", x"FF31", x"FF47", x"FF63", x"FF7C", x"FF99", x"FFA5", x"FFB6", x"FFB0", x"FFA7", x"FF91", x"FF77", x"FF5C", x"FF48", x"FF3C", x"FF38", x"FF36", x"FF3A", x"FF34", x"FF2F", x"FF28", x"FF28", x"FF22", x"FF22", x"FF24", x"FF26", x"FF2D", x"FF37", x"FF48", x"FF49", x"FF4B", x"FF40", x"FF32", x"FF1D", x"FF0E", x"FF00", x"FEEE", x"FEEE", x"FEE5", x"FEE8", x"FEE8", x"FEE5", x"FEE2", x"FEDB", x"FEDA", x"FED4", x"FED9", x"FED9", x"FEE1", x"FEE4", x"FEE7", x"FEED", x"FEE9", x"FEE9", x"FEE3", x"FECF", x"FEC8", x"FEB1", x"FEAD", x"FEAC", x"FEB8", x"FECB", x"FED7", x"FEEE", x"FEF7", x"FF00", x"FF04", x"FF0D", x"FF07", x"FF0B", x"FF08", x"FF0D", x"FF15", x"FF1E", x"FF2D", x"FF2F", x"FF36", x"FF2E", x"FF24", x"FF16", x"FF05", x"FEFE", x"FEF0", x"FEF3", x"FEF0", x"FEF1", x"FEEE", x"FEEB", x"FEE4", x"FEE2", x"FEDA", x"FED4", x"FED5", x"FECC", x"FED3", x"FED7", x"FEE1", x"FEEA", x"FEEE", x"FEED", x"FEE9", x"FED1", x"FEC3", x"FEA7", x"FE91", x"FE8E", x"FE88", x"FE96", x"FE97", x"FEAA", x"FEAE", x"FEBA", x"FEC9", x"FED3", x"FEE1", x"FEF4", x"FF07", x"FF1F", x"FF3F", x"FF64", x"FF81", x"FF97", x"FFA5", x"FFA3", x"FF9E", x"FF90", x"FF8A", x"FF7B", x"FF75", x"FF70", x"FF61", x"FF59", x"FF43", x"FF37", x"FF1A", x"FF0F", x"FEFB", x"FEF2", x"FEEC", x"FEEC", x"FEEE", x"FEF5", x"FEFC", x"FF07", x"FF0B", x"FF11", x"FF07", x"FEFB", x"FEE8", x"FED8", x"FECC", x"FECD", x"FED1", x"FED4", x"FEE0", x"FEDE", x"FEDD", x"FEDA", x"FEDE", x"FEDD", x"FEE4", x"FEE7", x"FEF6", x"FEFD", x"FF17", x"FF28", x"FF37", x"FF3D", x"FF38", x"FF2B", x"FF13", x"FEFE", x"FEE8", x"FECD", x"FEBE", x"FEB1", x"FEA7", x"FEA2", x"FEA3", x"FE9D", x"FEA6", x"FEAA", x"FEB8", x"FEC3", x"FED7", x"FEE6", x"FF03", x"FF16", x"FF31", x"FF43", x"FF4F", x"FF57", x"FF47", x"FF3C", x"FF21", x"FF05", x"FEF2", x"FEE9", x"FEE8", x"FEF1", x"FEFC", x"FF03", x"FF0A", x"FF10", x"FF1A", x"FF1C", x"FF2D", x"FF35", x"FF3E", x"FF4D", x"FF61", x"FF71", x"FF7F", x"FF88", x"FF7D", x"FF6F", x"FF50", x"FF3D", x"FF24", x"FF12", x"FF0B", x"FF03", x"FEF9", x"FEFF", x"FEF3", x"FEF9", x"FEF4", x"FEFB", x"FEF5", x"FF01", x"FF02", x"FF18", x"FF1B", x"FF35", x"FF41", x"FF53", x"FF5C", x"FF61", x"FF57", x"FF49", x"FF38", x"FF27", x"FF23", x"FF26", x"FF2F", x"FF41", x"FF48", x"FF59", x"FF5C", x"FF69", x"FF6A", x"FF75", x"FF78", x"FF84", x"FF8C", x"FF9F", x"FFAF", x"FFC0", x"FFCC", x"FFD0", x"FFCB", x"FFC0", x"FFAE", x"FFA2", x"FF93", x"FF8C", x"FF8B", x"FF80", x"FF81", x"FF77", x"FF71", x"FF67", x"FF5E", x"FF57", x"FF4E", x"FF4D", x"FF48", x"FF4D", x"FF52", x"FF5E", x"FF6B", x"FF7C", x"FF84", x"FF8A", x"FF81", x"FF74", x"FF62", x"FF57", x"FF4B", x"FF4F", x"FF51", x"FF61", x"FF69", x"FF6F", x"FF73", x"FF7B", x"FF7B", x"FF88", x"FF8F", x"FF9C", x"FFA4", x"FFC1", x"FFD7", x"FFF3", x"0011", x"0020", x"002C", x"0025", x"0025", x"001A", x"000D", x"0005", x"FFF7", x"FFE4", x"FFD7", x"FFCA", x"FFB1", x"FF9E", x"FF85", x"FF76", x"FF61", x"FF5F", x"FF57", x"FF5C", x"FF60", x"FF6E", x"FF79", x"FF8C", x"FF96", x"FF99", x"FF96", x"FF87", x"FF7A", x"FF68", x"FF66", x"FF65", x"FF74", x"FF77", x"FF8C", x"FF83", x"FF8D", x"FF8C", x"FF8C", x"FF92", x"FF9B", x"FF9D", x"FFB5", x"FFC4", x"FFE2", x"FFF2", x"000A", x"000F", x"0010", x"0008", x"FFFF", x"FFF5", x"FFE9", x"FFEC", x"FFE2", x"FFE5", x"FFE6", x"FFE4", x"FFE5", x"FFE5", x"FFE3", x"FFEB", x"FFEE", x"FFFD", x"000A", x"001D", x"0036", x"004C", x"0065", x"0079", x"0082", x"0081", x"007B", x"0068", x"0054", x"0044", x"0035", x"0034", x"0034", x"0040", x"003C", x"003E", x"003C", x"0037", x"003A", x"003D", x"003D", x"003C", x"0042", x"0053", x"005A", x"0071", x"007B", x"007A", x"0071", x"0068", x"005C", x"004E", x"0047", x"003E", x"0031", x"002A", x"002A", x"0023", x"0022", x"0025", x"0023", x"0027", x"0029", x"0032", x"0032", x"0033", x"003A", x"003B", x"0042", x"0043", x"0042", x"0030", x"0022", x"000C", x"FFFF", x"FFF7", x"FFFA", x"0006", x"001B", x"0030", x"0043", x"0053", x"005A", x"0060", x"0065", x"006A", x"006F", x"006F", x"007E", x"0083", x"0094", x"009D", x"00AA", x"009D", x"009D", x"008C", x"0082", x"0070", x"006B", x"005D", x"0059", x"0052", x"0053", x"0047", x"0042", x"0037", x"002E", x"0024", x"0020", x"001C", x"001B", x"001A", x"0022", x"0024", x"0034", x"0033", x"003C", x"0033", x"002B", x"001C", x"000E", x"0009", x"000A", x"0013", x"0027", x"0030", x"0041", x"0048", x"0058", x"005C", x"0074", x"007B", x"008F", x"009C", x"00B4", x"00CF", x"00E3", x"0105", x"010C", x"0117", x"0117", x"0116", x"0111", x"010C", x"010D", x"0101", x"00FF", x"00F8", x"00F4", x"00E8", x"00E2", x"00D5", x"00C7", x"00BC", x"00B7", x"00AE", x"00AC", x"00AC", x"00AE", x"00B1", x"00B9", x"00B7", x"00BA", x"00AB", x"00A6", x"008A", x"0081", x"0077", x"0078", x"007D", x"008E", x"0092", x"009D", x"00A2", x"00A6", x"00AB", x"00B2", x"00B6", x"00BB", x"00C0", x"00D2", x"00DB", x"00F0", x"00F9", x"00FB", x"00F1", x"00E3", x"00D0", x"00BC", x"00AC", x"009F", x"008F", x"0085", x"0086", x"007A", x"007E", x"0078", x"0081", x"0082", x"008C", x"009B", x"00A3", x"00B5", x"00C3", x"00D4", x"00E4", x"00F4", x"00F7", x"00FB", x"00EA", x"00D8", x"00C2", x"00A9", x"009E", x"0093", x"0098", x"00A2", x"00A7", x"00B4", x"00B8", x"00BF", x"00C6", x"00D3", x"00DD", x"00E1", x"00F6", x"00FE", x"010F", x"0123", x"012B", x"0132", x"0127", x"0124", x"010F", x"0102", x"00F4", x"00E4", x"00D3", x"00CC", x"00C2", x"00C0", x"00B7", x"00B4", x"00B1", x"00AB", x"00B3", x"00B5", x"00BF", x"00C7", x"00CF", x"00DB", x"00E4", x"00F4", x"00F6", x"00FA", x"00F4", x"00DD", x"00D1", x"00B9", x"00B7", x"00B5", x"00C6", x"00D4", x"00E0", x"00F2", x"00F6", x"0101", x"0109", x"0117", x"0114", x"0122", x"0125", x"0134", x"0135", x"014A", x"0141", x"0140", x"012F", x"0122", x"0108", x"00FB", x"00E8", x"00DA", x"00CE", x"00C3", x"00C3", x"00B9", x"00B8", x"00B3", x"00B0", x"00AC", x"00B8", x"00B3", x"00C4", x"00C8", x"00D5", x"00DB", x"00E9", x"00F0", x"00F8", x"00F1", x"00E8", x"00D2", x"00BE", x"00B0", x"00A1", x"00A4", x"00A7", x"00AE", x"00B8", x"00BF", x"00C6", x"00CB", x"00D7", x"00DC", x"00E8", x"00F5", x"0105", x"011A", x"0134", x"014D", x"0160", x"016B", x"0174", x"016B", x"0164", x"015A", x"014D", x"013D", x"012A", x"011B", x"0100", x"00F1", x"00DF", x"00D0", x"00C0", x"00B2", x"00AE", x"00A1", x"00A6", x"00A1", x"00A7", x"00AA", x"00B2", x"00BD", x"00BE", x"00C4", x"00B6", x"00A4", x"0094", x"0082", x"007A", x"007E", x"0083", x"0088", x"008C", x"008F", x"008F", x"0090", x"0097", x"0097", x"0097", x"00A3", x"00A8", x"00BC", x"00C9", x"00DC", x"00E3", x"00E3", x"00E1", x"00DA", x"00CD", x"00C8", x"00BF", x"00B4", x"00B2", x"00B2", x"00AF", x"00B2", x"00B0", x"00B1", x"00B0", x"00B8", x"00BC", x"00C7", x"00CD", x"00DD", x"00E5", x"00F4", x"0101", x"0107", x"010B", x"0104", x"00F5", x"00DB", x"00C7", x"00AB", x"009F", x"0098", x"0097", x"0094", x"0091", x"0091", x"0084", x"0087", x"0084", x"0081", x"0085", x"0088", x"0095", x"00A0", x"00B2", x"00C0", x"00C4", x"00CB", x"00C4", x"00BE", x"00AF", x"00A2", x"0095", x"0080", x"0077", x"0067", x"005E", x"0057", x"0052", x"0050", x"0052", x"0056", x"005A", x"005D", x"0064", x"0067", x"006A", x"0073", x"0072", x"0078", x"0077", x"006D", x"0062", x"004E", x"0042", x"0034", x"0037", x"003E", x"004A", x"0052", x"005E", x"005D", x"0060", x"0061", x"0061", x"005B", x"005A", x"005B", x"0054", x"0065", x"0068", x"0074", x"0070", x"0070", x"0063", x"0054", x"004D", x"0043", x"0036", x"002C", x"0026", x"001C", x"0016", x"0015", x"000E", x"0003", x"FFFE", x"FFF3", x"FFF0", x"FFEB", x"FFEF", x"FFEA", x"FFEB", x"FFF2", x"FFF7", x"FFF9", x"FFFD", x"FFF0", x"FFE4", x"FFCE", x"FFC3", x"FFB5", x"FFBB", x"FFBF", x"FFD0", x"FFDE", x"FFEB", x"FFFC", x"000A", x"0014", x"0025", x"002A", x"003B", x"0041", x"0055", x"0065", x"007B", x"0085", x"0092", x"0090", x"008F", x"0085", x"007E", x"006C", x"0064", x"0051", x"0047", x"0037", x"002C", x"0024", x"0017", x"0013", x"000B", x"0006", x"0001", x"FFFF", x"0000", x"FFFC", x"0001", x"0002", x"0001", x"0006", x"0004", x"FFF7", x"FFE9", x"FFD4", x"FFC3", x"FFB5", x"FFB6", x"FFB6", x"FFBD", x"FFBA", x"FFBF", x"FFB6", x"FFB6", x"FFB5", x"FFB3", x"FFB3", x"FFB3", x"FFB8", x"FFBE", x"FFC7", x"FFD6", x"FFD9", x"FFE0", x"FFDB", x"FFD4", x"FFC4", x"FFB9", x"FFA4", x"FF98", x"FF89", x"FF79", x"FF70", x"FF6D", x"FF68", x"FF67", x"FF68", x"FF6A", x"FF6B", x"FF79", x"FF7E", x"FF8B", x"FF8E", x"FF99", x"FFA0", x"FFA0", x"FFAB", x"FFA1", x"FF98", x"FF7F", x"FF71", x"FF59", x"FF57", x"FF52", x"FF5B", x"FF57", x"FF65", x"FF68", x"FF70", x"FF7A", x"FF80", x"FF82", x"FF88", x"FF8A", x"FF90", x"FF95", x"FFA0", x"FFA5", x"FFA9", x"FFAD", x"FFA0", x"FF99", x"FF84", x"FF7A", x"FF65", x"FF57", x"FF4B", x"FF3F", x"FF37", x"FF37", x"FF30", x"FF34", x"FF32", x"FF37", x"FF3D", x"FF42", x"FF4D", x"FF4E", x"FF57", x"FF5A", x"FF61", x"FF63", x"FF68", x"FF5F", x"FF50", x"FF44", x"FF31", x"FF29", x"FF20", x"FF2C", x"FF2E", x"FF3B", x"FF46", x"FF4D", x"FF57", x"FF60", x"FF67", x"FF71", x"FF78", x"FF80", x"FF88", x"FF91", x"FFA5", x"FFA8", x"FFB1", x"FFAD", x"FF9C", x"FF8D", x"FF79", x"FF66", x"FF50", x"FF3F", x"FF2C", x"FF1E", x"FF0F", x"FF08", x"FEFC", x"FEF0", x"FEF3", x"FEE7", x"FEF3", x"FEF9", x"FF07", x"FF0B", x"FF1B", x"FF1F", x"FF2C", x"FF2F", x"FF38", x"FF30", x"FF28", x"FF1A", x"FF0A", x"FF03", x"FEFE", x"FF05", x"FF0C", x"FF11", x"FF21", x"FF1F", x"FF2D", x"FF32", x"FF37", x"FF3C", x"FF42", x"FF46", x"FF54", x"FF5F", x"FF71", x"FF80", x"FF8A", x"FF94", x"FF91", x"FF8D", x"FF7F", x"FF70", x"FF5D", x"FF47", x"FF33", x"FF1B", x"FF10", x"FEFB", x"FEF3", x"FEE6", x"FEE1", x"FED7", x"FED8", x"FEDD", x"FED8", x"FEDF", x"FEE2", x"FEEC", x"FEF4", x"FF00", x"FF05", x"FEFE", x"FEF6", x"FEE2", x"FED4", x"FEC5", x"FEBE", x"FEC2", x"FEBF", x"FECB", x"FED2", x"FED7", x"FEE1", x"FEEA", x"FEED", x"FEF8", x"FF02", x"FF0F", x"FF20", x"FF2F", x"FF40", x"FF4E", x"FF54", x"FF5B", x"FF54", x"FF4E", x"FF45", x"FF37", x"FF2C", x"FF21", x"FF19", x"FF11", x"FF10", x"FF0B", x"FF0C", x"FF0C", x"FF0D", x"FF15", x"FF1D", x"FF2E", x"FF3B", x"FF47", x"FF59", x"FF5D", x"FF6C", x"FF6F", x"FF6C", x"FF62", x"FF53", x"FF3D", x"FF2B", x"FF1A", x"FF13", x"FF0E", x"FF05", x"FF0E", x"FF07", x"FF0D", x"FF13", x"FF18", x"FF1A", x"FF1D", x"FF1D", x"FF25", x"FF2A", x"FF3E", x"FF49", x"FF59", x"FF63", x"FF6C", x"FF6E", x"FF6C", x"FF67", x"FF57", x"FF49", x"FF3A", x"FF27", x"FF1F", x"FF11", x"FF09", x"FF06", x"FF05", x"FF04", x"FF0D", x"FF0C", x"FF1A", x"FF13", x"FF20", x"FF17", x"FF1D", x"FF1D", x"FF22", x"FF21", x"FF19", x"FF13", x"FEFF", x"FEF8", x"FEF5", x"FEF9", x"FF00", x"FF0C", x"FF1A", x"FF24", x"FF30", x"FF3D", x"FF45", x"FF45", x"FF4B", x"FF4C", x"FF4E", x"FF5C", x"FF60", x"FF6C", x"FF69", x"FF6F", x"FF65", x"FF5C", x"FF4B", x"FF3C", x"FF2A", x"FF1B", x"FF13", x"FF04", x"FEFD", x"FEF6", x"FEEA", x"FEE9", x"FEE3", x"FEDD", x"FEE3", x"FEE2", x"FEEC", x"FEF0", x"FEFA", x"FF02", x"FF06", x"FF11", x"FF18", x"FF1C", x"FF14", x"FF0F", x"FEFA", x"FEF8", x"FEED", x"FEF8", x"FEFB", x"FF0B", x"FF1A", x"FF28", x"FF37", x"FF47", x"FF52", x"FF5D", x"FF6C", x"FF78", x"FF87", x"FF9B", x"FFAC", x"FFBF", x"FFD0", x"FFDF", x"FFE3", x"FFED", x"FFE7", x"FFE4", x"FFD7", x"FFD2", x"FFB8", x"FFB4", x"FF9F", x"FF98", x"FF8D", x"FF8D", x"FF87", x"FF89", x"FF87", x"FF8C", x"FF89", x"FF8D", x"FF8B", x"FF8F", x"FF94", x"FFA1", x"FFA2", x"FFA5", x"FF9A", x"FF94", x"FF7F", x"FF79", x"FF72", x"FF71", x"FF73", x"FF79", x"FF80", x"FF87", x"FF8D", x"FF92", x"FF91", x"FF9A", x"FF9B", x"FFA4", x"FFAC", x"FFBC", x"FFCA", x"FFD3", x"FFE2", x"FFE7", x"FFE8", x"FFE7", x"FFE3", x"FFD3", x"FFCC", x"FFBC", x"FFAF", x"FFA8", x"FFA0", x"FFA2", x"FFA0", x"FFA8", x"FFA9", x"FFB5", x"FFB8", x"FFC4", x"FFC6", x"FFD0", x"FFD2", x"FFD7", x"FFDB", x"FFDA", x"FFDA", x"FFC8", x"FFBD", x"FFA2", x"FF8E", x"FF83", x"FF7C", x"FF78", x"FF7C", x"FF81", x"FF85", x"FF94", x"FFA2", x"FFB4", x"FFC2", x"FFCC", x"FFDC", x"FFDE", x"FFF4", x"FFFF", x"0015", x"001F", x"002E", x"0032", x"0035", x"0030", x"0026", x"0018", x"0006", x"FFF4", x"FFE4", x"FFD8", x"FFCA", x"FFC6", x"FFC2", x"FFC4", x"FFC9", x"FFD5", x"FFDB", x"FFEC", x"FFEE", x"FFFE", x"0004", x"000A", x"001B", x"001D", x"0022", x"0020", x"001A", x"0010", x"0002", x"0006", x"FFFF", x"000C", x"0016", x"001E", x"002B", x"0031", x"0043", x"004A", x"005A", x"0063", x"006B", x"0070", x"0078", x"0082", x"0088", x"008E", x"008E", x"0087", x"0080", x"0076", x"0067", x"0058", x"004B", x"0038", x"002C", x"0021", x"0020", x"001A", x"0020", x"0024", x"0029", x"0032", x"003D", x"0043", x"004B", x"0053", x"0052", x"005D", x"005A", x"0063", x"005C", x"0057", x"004B", x"003D", x"0031", x"002D", x"002E", x"0033", x"0040", x"004D", x"0059", x"0068", x"0076", x"007E", x"008A", x"008F", x"0093", x"009C", x"00A8", x"00B3", x"00C5", x"00CE", x"00DC", x"00DE", x"00E4", x"00E2", x"00D6", x"00CD", x"00B7", x"00A3", x"0090", x"007E", x"0072", x"0064", x"0062", x"0057", x"005E", x"0057", x"005D", x"005E", x"0062", x"006E", x"0072", x"007F", x"008B", x"008A", x"0094", x"0089", x"0081", x"0070", x"0063", x"005A", x"004F", x"0054", x"004C", x"004F", x"0049", x"0053", x"0057", x"0063", x"0070", x"007B", x"0083", x"0094", x"009C", x"00B0", x"00B8", x"00C9", x"00CA", x"00D3", x"00D3", x"00D4", x"00D0", x"00C9", x"00BF", x"00B3", x"00AB", x"00A6", x"009E", x"00A4", x"00A4", x"00A7", x"00AB", x"00B5", x"00B9", x"00C2", x"00CA", x"00D1", x"00D7", x"00DF", x"00EA", x"00E7", x"00E9", x"00DC", x"00D2", x"00BE", x"00B4", x"00AA", x"00A0", x"009D", x"009A", x"0096", x"009B", x"00A2", x"00A9", x"00B6", x"00BA", x"00C4", x"00C8", x"00D3", x"00DA", x"00E5", x"00F3", x"0104", x"010E", x"011A", x"011A", x"0115", x"0109", x"00FA", x"00E2", x"00D2", x"00BA", x"00AF", x"00A3", x"00A2", x"00A0", x"00A2", x"00A5", x"00B4", x"00B7", x"00CA", x"00D2", x"00DD", x"00E7", x"00EC", x"00F1", x"00F4", x"00EE", x"00E7", x"00D9", x"00CE", x"00C6", x"00BD", x"00BF", x"00C0", x"00C0", x"00C4", x"00C6", x"00D5", x"00D7", x"00E9", x"00EA", x"00F2", x"00F7", x"00FF", x"0104", x"010A", x"0112", x"0110", x"010F", x"0107", x"0102", x"00F7", x"00EB", x"00DE", x"00CE", x"00BA", x"00B4", x"00A5", x"00A4", x"00A4", x"00A3", x"00A8", x"00AB", x"00AC", x"00AF", x"00B7", x"00B8", x"00C4", x"00C4", x"00CE", x"00D2", x"00CF", x"00D1", x"00CA", x"00C1", x"00BA", x"00B5", x"00B2", x"00B8", x"00BD", x"00C6", x"00CE", x"00E2", x"00ED", x"0101", x"010B", x"0116", x"0117", x"011C", x"0122", x"012A", x"0136", x"0145", x"014D", x"015A", x"015F", x"0160", x"0161", x"0154", x"014E", x"013A", x"012C", x"0119", x"010A", x"0102", x"00F9", x"00FA", x"00F4", x"00FD", x"00F9", x"00FE", x"00FE", x"0100", x"00FD", x"0100", x"0101", x"00FE", x"00F7", x"00EF", x"00DA", x"00D0", x"00BC", x"00B8", x"00AB", x"00AA", x"00A3", x"00A2", x"009C", x"00A0", x"00A0", x"00A3", x"00A8", x"00A8", x"00AD", x"00AD", x"00B2", x"00B7", x"00C7", x"00CE", x"00DA", x"00E1", x"00E7", x"00E6", x"00E5", x"00D9", x"00D0", x"00BC", x"00B4", x"00A6", x"00A1", x"009E", x"009C", x"009B", x"009E", x"00A0", x"00A4", x"00A9", x"00AA", x"00B3", x"00B2", x"00C0", x"00C0", x"00C7", x"00C5", x"00BD", x"00B7", x"00A6", x"00A3", x"0096", x"0090", x"0091", x"008A", x"008B", x"008D", x"0091", x"0098", x"009D", x"00A5", x"00A4", x"00A7", x"00AA", x"00AC", x"00B6", x"00C1", x"00C9", x"00CF", x"00D0", x"00D1", x"00C8", x"00C3", x"00B3", x"00A2", x"008C", x"007D", x"006B", x"005F", x"0059", x"0052", x"0051", x"0054", x"004D", x"0057", x"0053", x"0060", x"0063", x"006F", x"0076", x"007A", x"007C", x"007A", x"006F", x"0069", x"0060", x"005F", x"0056", x"005A", x"0058", x"005A", x"005B", x"0065", x"006F", x"007D", x"008C", x"0094", x"009B", x"00A2", x"00A5", x"00B0", x"00AD", x"00B9", x"00B8", x"00B9", x"00AF", x"00A6", x"0094", x"0080", x"006E", x"0057", x"0045", x"0037", x"0026", x"0028", x"0020", x"002A", x"002D", x"0035", x"0037", x"003D", x"003F", x"0045", x"0047", x"004D", x"0053", x"0052", x"0054", x"0051", x"0042", x"003B", x"0027", x"0028", x"001A", x"0022", x"001B", x"0021", x"0026", x"002C", x"003A", x"0041", x"0049", x"0050", x"004F", x"0051", x"0058", x"0053", x"0060", x"005F", x"0069", x"006B", x"006F", x"0069", x"0060", x"0055", x"0044", x"0032", x"0024", x"0010", x"FFFF", x"FFF1", x"FFE2", x"FFDC", x"FFD1", x"FFD0", x"FFCA", x"FFC8", x"FFC7", x"FFC5", x"FFC5", x"FFC8", x"FFC5", x"FFCA", x"FFC1", x"FFBD", x"FFB6", x"FFA8", x"FFA6", x"FFA0", x"FF9D", x"FFA0", x"FF98", x"FF9C", x"FF9D", x"FFA3", x"FFAE", x"FFB8", x"FFC7", x"FFD0", x"FFDA", x"FFE0", x"FFE8", x"FFEE", x"FFF3", x"FFF8", x"FFF8", x"FFFD", x"FFFA", x"FFFA", x"FFF4", x"FFEF", x"FFE9", x"FFE1", x"FFDA", x"FFDB", x"FFD3", x"FFD6", x"FFD3", x"FFD9", x"FFD4", x"FFDE", x"FFD4", x"FFE0", x"FFDA", x"FFE1", x"FFE5", x"FFE8", x"FFEA", x"FFE9", x"FFE1", x"FFDA", x"FFC7", x"FFBD", x"FFB0", x"FFA8", x"FFA6", x"FFA1", x"FF9E", x"FF97", x"FF98", x"FF9F", x"FFA1", x"FFAF", x"FFB2", x"FFB8", x"FFC0", x"FFC7", x"FFD4", x"FFDD", x"FFF1", x"FFFF", x"000B", x"0014", x"0017", x"0015", x"0006", x"FFFF", x"FFE8", x"FFDB", x"FFBF", x"FFAF", x"FF97", x"FF89", x"FF7B", x"FF76", x"FF70", x"FF6E", x"FF6C", x"FF6F", x"FF74", x"FF7F", x"FF87", x"FF91", x"FF94", x"FF93", x"FF8C", x"FF81", x"FF74", x"FF69", x"FF63", x"FF5D", x"FF5A", x"FF5B", x"FF53", x"FF56", x"FF54", x"FF5B", x"FF60", x"FF6B", x"FF71", x"FF74", x"FF78", x"FF73", x"FF79", x"FF70", x"FF7B", x"FF71", x"FF77", x"FF6A", x"FF66", x"FF55", x"FF48", x"FF32", x"FF22", x"FF0F", x"FF05", x"FEF9", x"FEF4", x"FEF2", x"FEF2", x"FEF5", x"FEF9", x"FEFA", x"FF00", x"FEFE", x"FF03", x"FF0A", x"FF0E", x"FF1B", x"FF20", x"FF22", x"FF21", x"FF18", x"FF15", x"FF08", x"FF06", x"FF00", x"FEFD", x"FEFD", x"FEFF", x"FF02", x"FF13", x"FF1C", x"FF32", x"FF3E", x"FF50", x"FF50", x"FF60", x"FF5E", x"FF6C", x"FF70", x"FF80", x"FF84", x"FF92", x"FF96", x"FF98", x"FF94", x"FF8A", x"FF7E", x"FF71", x"FF62", x"FF52", x"FF46", x"FF33", x"FF31", x"FF2A", x"FF2B", x"FF30", x"FF32", x"FF36", x"FF39", x"FF3C", x"FF43", x"FF43", x"FF48", x"FF42", x"FF3D", x"FF31", x"FF23", x"FF18", x"FF0B", x"FF03", x"FEFB", x"FEF7", x"FEEB", x"FEE7", x"FEE1", x"FEE1", x"FEEA", x"FEEF", x"FF00", x"FF06", x"FF0C", x"FF13", x"FF18", x"FF1C", x"FF23", x"FF2A", x"FF32", x"FF3C", x"FF3E", x"FF44", x"FF41", x"FF42", x"FF43", x"FF41", x"FF41", x"FF40", x"FF38", x"FF37", x"FF2F", x"FF31", x"FF2A", x"FF27", x"FF1F", x"FF1A", x"FF16", x"FF13", x"FF17", x"FF19", x"FF1F", x"FF1A", x"FF21", x"FF12", x"FF10", x"FF01", x"FEFF", x"FEFA", x"FEF4", x"FEFA", x"FEEE", x"FEEF", x"FEED", x"FEF3", x"FEFA", x"FF04", x"FF0F", x"FF16", x"FF1C", x"FF26", x"FF2D", x"FF39", x"FF44", x"FF4F", x"FF52", x"FF5C", x"FF56", x"FF55", x"FF47", x"FF3F", x"FF33", x"FF22", x"FF17", x"FF0E", x"FEFE", x"FEFC", x"FEF4", x"FEEE", x"FEEF", x"FEE8", x"FEE9", x"FEE9", x"FEEF", x"FEFF", x"FF08", x"FF1F", x"FF28", x"FF35", x"FF39", x"FF36", x"FF35", x"FF2E", x"FF2C", x"FF29", x"FF2B", x"FF2B", x"FF2B", x"FF2B", x"FF2D", x"FF32", x"FF34", x"FF42", x"FF44", x"FF4C", x"FF54", x"FF53", x"FF5B", x"FF5C", x"FF65", x"FF6A", x"FF70", x"FF6D", x"FF64", x"FF5A", x"FF47", x"FF3B", x"FF2C", x"FF1E", x"FF1C", x"FF0E", x"FF12", x"FF0E", x"FF12", x"FF15", x"FF14", x"FF16", x"FF12", x"FF13", x"FF13", x"FF1B", x"FF23", x"FF27", x"FF33", x"FF2F", x"FF34", x"FF2C", x"FF28", x"FF23", x"FF18", x"FF1D", x"FF19", x"FF1E", x"FF20", x"FF2B", x"FF32", x"FF42", x"FF50", x"FF5F", x"FF69", x"FF6E", x"FF72", x"FF77", x"FF75", x"FF7E", x"FF82", x"FF86", x"FF91", x"FF90", x"FF91", x"FF86", x"FF7F", x"FF74", x"FF6A", x"FF66", x"FF59", x"FF55", x"FF45", x"FF48", x"FF3C", x"FF45", x"FF40", x"FF49", x"FF47", x"FF4C", x"FF4B", x"FF56", x"FF5B", x"FF61", x"FF67", x"FF63", x"FF5E", x"FF53", x"FF46", x"FF3D", x"FF37", x"FF32", x"FF2F", x"FF2E", x"FF2B", x"FF29", x"FF2E", x"FF33", x"FF41", x"FF4E", x"FF5B", x"FF64", x"FF6D", x"FF73", x"FF78", x"FF82", x"FF86", x"FF91", x"FF93", x"FF96", x"FF92", x"FF8E", x"FF8B", x"FF86", x"FF8A", x"FF87", x"FF87", x"FF86", x"FF86", x"FF82", x"FF87", x"FF7B", x"FF7E", x"FF75", x"FF78", x"FF76", x"FF78", x"FF82", x"FF84", x"FF8B", x"FF91", x"FF8D", x"FF89", x"FF7E", x"FF7B", x"FF6E", x"FF72", x"FF6F", x"FF79", x"FF76", x"FF7D", x"FF7E", x"FF83", x"FF8B", x"FF97", x"FF9D", x"FFA9", x"FFB1", x"FFB9", x"FFBF", x"FFC8", x"FFD4", x"FFDA", x"FFE5", x"FFE6", x"FFE5", x"FFE3", x"FFD9", x"FFD6", x"FFCA", x"FFC6", x"FFBF", x"FFBA", x"FFB4", x"FFB0", x"FFAF", x"FFAA", x"FFAC", x"FFA7", x"FFB1", x"FFAF", x"FFBD", x"FFC6", x"FFD4", x"FFE0", x"FFEB", x"FFF2", x"FFF1", x"FFF0", x"FFE3", x"FFDC", x"FFCC", x"FFC8", x"FFBE", x"FFBE", x"FFB7", x"FFBC", x"FFB1", x"FFB9", x"FFBB", x"FFC4", x"FFCA", x"FFD6", x"FFDC", x"FFDF", x"FFE6", x"FFE7", x"FFEA", x"FFF4", x"FFEC", x"FFF5", x"FFDE", x"FFDA", x"FFC3", x"FFB3", x"FFA9", x"FF9C", x"FF9C", x"FF94", x"FF99", x"FF95", x"FF9F", x"FFA2", x"FFA6", x"FFAC", x"FFAD", x"FFB1", x"FFBA", x"FFC2", x"FFD1", x"FFD8", x"FFE4", x"FFEE", x"FFF1", x"FFF7", x"FFF5", x"FFEC", x"FFED", x"FFE6", x"FFEC", x"FFE8", x"FFEE", x"FFED", x"FFF3", x"FFFA", x"0008", x"0011", x"0022", x"002B", x"0034", x"003B", x"0041", x"004F", x"0054", x"0065", x"006B", x"0076", x"0070", x"0072", x"0065", x"0065", x"0059", x"005A", x"004D", x"004D", x"0040", x"0044", x"003F", x"0043", x"0045", x"0047", x"004B", x"004C", x"0056", x"005A", x"005D", x"0061", x"0061", x"0061", x"0057", x"0054", x"0040", x"0039", x"002C", x"0026", x"001E", x"001B", x"0015", x"0013", x"0013", x"0019", x"001E", x"002A", x"0038", x"0047", x"0051", x"005D", x"0065", x"0069", x"0076", x"007A", x"0084", x"0085", x"0087", x"0083", x"0080", x"007C", x"007D", x"0073", x"0077", x"0071", x"006E", x"006A", x"0069", x"005C", x"005C", x"004F", x"0052", x"004B", x"0051", x"0054", x"0058", x"0063", x"0069", x"0070", x"0070", x"0071", x"006F", x"0068", x"0066", x"0061", x"005C", x"0061", x"005A", x"005A", x"0055", x"0059", x"0057", x"0060", x"006B", x"006F", x"007E", x"007F", x"008D", x"0094", x"00A1", x"00A9", x"00B0", x"00AF", x"00AD", x"00A3", x"00A0", x"0093", x"0092", x"0087", x"0087", x"007E", x"0075", x"0074", x"0069", x"0066", x"0069", x"0060", x"0069", x"0065", x"0073", x"007A", x"0086", x"0092", x"009B", x"009D", x"00A5", x"009C", x"009C", x"0093", x"0090", x"0092", x"0092", x"009C", x"009B", x"009F", x"00A6", x"00A5", x"00B2", x"00B3", x"00C2", x"00C1", x"00CC", x"00D0", x"00D4", x"00DE", x"00E0", x"00E5", x"00E3", x"00DE", x"00D1", x"00C8", x"00B9", x"00B3", x"00AC", x"00A8", x"00A9", x"00A2", x"00AA", x"00A5", x"00AA", x"00A7", x"00AA", x"00A8", x"00A9", x"00AE", x"00B7", x"00BB", x"00C4", x"00CB", x"00CF", x"00D3", x"00D0", x"00CD", x"00C4", x"00C0", x"00BC", x"00B7", x"00BB", x"00BA", x"00BF", x"00C2", x"00C5", x"00CD", x"00D0", x"00DD", x"00DE", x"00EA", x"00EB", x"00F3", x"00F5", x"00FD", x"0105", x"010B", x"0111", x"010B", x"010C", x"0100", x"0101", x"00F6", x"00F7", x"00ED", x"00EE", x"00E3", x"00E6", x"00DE", x"00E0", x"00D6", x"00D6", x"00CF", x"00CB", x"00CE", x"00C3", x"00CF", x"00C6", x"00D3", x"00CD", x"00D0", x"00C8", x"00C4", x"00BB", x"00B7", x"00B5", x"00B7", x"00B9", x"00C3", x"00C2", x"00CD", x"00C9", x"00CF", x"00D0", x"00D7", x"00DC", x"00E2", x"00E7", x"00E9", x"00EB", x"00F4", x"00F9", x"00FC", x"0100", x"00FA", x"00FB", x"00F2", x"00F9", x"00F3", x"00FA", x"00FD", x"00FE", x"0100", x"0101", x"00FD", x"00FB", x"00F3", x"00EF", x"00E3", x"00E5", x"00DB", x"00E1", x"00DE", x"00E6", x"00E4", x"00E6", x"00E4", x"00E2", x"00D6", x"00D2", x"00C9", x"00C1", x"00C6", x"00C1", x"00C9", x"00C4", x"00C9", x"00C9", x"00D1", x"00D6", x"00E4", x"00E9", x"00F7", x"00FB", x"0108", x"010E", x"0115", x"011A", x"011D", x"011A", x"0113", x"0106", x"00FB", x"00EC", x"00E5", x"00DE", x"00D3", x"00CA", x"00BA", x"00B6", x"00A8", x"00A9", x"00A0", x"00A3", x"009E", x"00A5", x"00A7", x"00AF", x"00B7", x"00C4", x"00C7", x"00D5", x"00D3", x"00D0", x"00C5", x"00B9", x"00AE", x"00A6", x"00A1", x"009D", x"0096", x"0093", x"008E", x"008A", x"008E", x"008C", x"0096", x"0097", x"009E", x"009F", x"00A0", x"00A4", x"00A5", x"00A4", x"00A3", x"0094", x"0083", x"0073", x"005F", x"0057", x"0048", x"004A", x"003F", x"0044", x"0040", x"0049", x"0046", x"004D", x"004A", x"004A", x"004C", x"004E", x"0054", x"0055", x"005D", x"0060", x"0064", x"0068", x"0064", x"0066", x"0053", x"005A", x"0046", x"0052", x"004E", x"0055", x"005B", x"005B", x"0065", x"0063", x"006B", x"0071", x"0079", x"0081", x"0088", x"008C", x"008E", x"0094", x"0092", x"0099", x"0095", x"0091", x"008B", x"007E", x"007D", x"006E", x"006E", x"0066", x"0061", x"005F", x"0056", x"0056", x"004F", x"0052", x"004C", x"004E", x"004C", x"004D", x"004E", x"0051", x"0055", x"0052", x"0052", x"004C", x"0042", x"0038", x"0026", x"001D", x"000A", x"0006", x"0000", x"FFFF", x"0001", x"FFFE", x"FFFD", x"FFFE", x"0000", x"000B", x"000F", x"001D", x"0025", x"002F", x"003A", x"0041", x"004D", x"0052", x"005C", x"0058", x"0057", x"0052", x"004D", x"004A", x"004E", x"004A", x"0049", x"0045", x"0039", x"0030", x"0025", x"0018", x"000B", x"FFFC", x"FFF1", x"FFEC", x"FFE4", x"FFE2", x"FFE7", x"FFE5", x"FFEE", x"FFEF", x"FFF2", x"FFEA", x"FFE5", x"FFDA", x"FFD8", x"FFD3", x"FFD8", x"FFD5", x"FFD9", x"FFD3", x"FFD5", x"FFCB", x"FFD3", x"FFC9", x"FFD6", x"FFD0", x"FFDE", x"FFDC", x"FFE4", x"FFEC", x"FFF0", x"FFF7", x"FFF8", x"FFF3", x"FFEB", x"FFE0", x"FFD6", x"FFCC", x"FFCA", x"FFBF", x"FFBA", x"FFB6", x"FFAF", x"FFAB", x"FFA4", x"FFA2", x"FF9D", x"FFA0", x"FFA6", x"FFAE", x"FFB7", x"FFC2", x"FFCC", x"FFD9", x"FFE3", x"FFE8", x"FFE8", x"FFE0", x"FFD2", x"FFCA", x"FFBD", x"FFBB", x"FFBA", x"FFB8", x"FFBB", x"FFB5", x"FFB6", x"FFB0", x"FFB3", x"FFB4", x"FFBE", x"FFC5", x"FFCC", x"FFD5", x"FFD8", x"FFE1", x"FFE3", x"FFE4", x"FFDD", x"FFD5", x"FFC7", x"FFBE", x"FFAF", x"FFAC", x"FFA7", x"FFA5", x"FFAB", x"FFA4", x"FFAB", x"FFA2", x"FFA3", x"FF9F", x"FF95", x"FF95", x"FF8D", x"FF91", x"FF8E", x"FF94", x"FF96", x"FF9C", x"FF9F", x"FFA5", x"FF99", x"FF9A", x"FF89", x"FF87", x"FF7B", x"FF81", x"FF82", x"FF86", x"FF8A", x"FF8A", x"FF88", x"FF8A", x"FF8E", x"FF8F", x"FF97", x"FF95", x"FF9F", x"FF99", x"FFA4", x"FF9F", x"FFA3", x"FF9E", x"FF9A", x"FF8F", x"FF89", x"FF7D", x"FF77", x"FF73", x"FF73", x"FF6F", x"FF75", x"FF6E", x"FF74", x"FF6B", x"FF6D", x"FF63", x"FF5C", x"FF57", x"FF4E", x"FF4D", x"FF47", x"FF4B", x"FF47", x"FF4C", x"FF45", x"FF46", x"FF3A", x"FF2F", x"FF26", x"FF17", x"FF1D", x"FF1B", x"FF29", x"FF2D", x"FF36", x"FF39", x"FF3C", x"FF3C", x"FF3E", x"FF3E", x"FF45", x"FF48", x"FF4F", x"FF57", x"FF5D", x"FF69", x"FF6A", x"FF71", x"FF6B", x"FF65", x"FF5C", x"FF55", x"FF4F", x"FF54", x"FF53", x"FF57", x"FF56", x"FF52", x"FF4C", x"FF40", x"FF39", x"FF2A", x"FF22", x"FF19", x"FF13", x"FF11", x"FF11", x"FF14", x"FF18", x"FF21", x"FF28", x"FF32", x"FF2B", x"FF2A", x"FF21", x"FF1B", x"FF22", x"FF25", x"FF2B", x"FF31", x"FF33", x"FF31", x"FF32", x"FF2E", x"FF32", x"FF33", x"FF3C", x"FF40", x"FF49", x"FF4C", x"FF55", x"FF58", x"FF5D", x"FF60", x"FF5B", x"FF5B", x"FF4F", x"FF49", x"FF44", x"FF41", x"FF41", x"FF40", x"FF40", x"FF3E", x"FF3C", x"FF34", x"FF33", x"FF2A", x"FF28", x"FF2A", x"FF2A", x"FF32", x"FF3C", x"FF46", x"FF51", x"FF59", x"FF5E", x"FF5A", x"FF4E", x"FF43", x"FF30", x"FF25", x"FF1D", x"FF17", x"FF13", x"FF17", x"FF12", x"FF15", x"FF11", x"FF10", x"FF13", x"FF11", x"FF1A", x"FF1C", x"FF23", x"FF2A", x"FF2A", x"FF34", x"FF2B", x"FF2C", x"FF1C", x"FF11", x"FF00", x"FEF5", x"FEE9", x"FEE6", x"FEE2", x"FEE7", x"FEE8", x"FEF0", x"FEEF", x"FEF7", x"FEF3", x"FEF9", x"FEF7", x"FF00", x"FEFE", x"FF08", x"FF0F", x"FF17", x"FF23", x"FF2B", x"FF35", x"FF2D", x"FF2C", x"FF20", x"FF17", x"FF15", x"FF19", x"FF20", x"FF2A", x"FF31", x"FF37", x"FF37", x"FF3C", x"FF42", x"FF42", x"FF4C", x"FF50", x"FF57", x"FF5E", x"FF61", x"FF67", x"FF6E", x"FF6A", x"FF6E", x"FF64", x"FF5C", x"FF59", x"FF4E", x"FF52", x"FF4F", x"FF53", x"FF56", x"FF57", x"FF59", x"FF56", x"FF55", x"FF4D", x"FF49", x"FF42", x"FF41", x"FF3C", x"FF42", x"FF3C", x"FF45", x"FF3F", x"FF47", x"FF41", x"FF40", x"FF37", x"FF29", x"FF1C", x"FF14", x"FF14", x"FF17", x"FF21", x"FF27", x"FF2F", x"FF31", x"FF39", x"FF39", x"FF41", x"FF46", x"FF4C", x"FF58", x"FF5B", x"FF67", x"FF6B", x"FF73", x"FF77", x"FF76", x"FF78", x"FF6F", x"FF73", x"FF69", x"FF71", x"FF72", x"FF75", x"FF7A", x"FF79", x"FF77", x"FF76", x"FF6C", x"FF65", x"FF58", x"FF52", x"FF47", x"FF48", x"FF48", x"FF4D", x"FF4D", x"FF58", x"FF5A", x"FF67", x"FF64", x"FF65", x"FF5F", x"FF54", x"FF57", x"FF55", x"FF5A", x"FF5D", x"FF63", x"FF5E", x"FF62", x"FF56", x"FF5A", x"FF54", x"FF58", x"FF5F", x"FF64", x"FF6D", x"FF76", x"FF7C", x"FF84", x"FF88", x"FF89", x"FF88", x"FF82", x"FF82", x"FF7A", x"FF7E", x"FF7B", x"FF7C", x"FF7C", x"FF79", x"FF79", x"FF75", x"FF71", x"FF6D", x"FF68", x"FF71", x"FF6D", x"FF80", x"FF88", x"FF96", x"FFA7", x"FFAA", x"FFB7", x"FFB1", x"FFB0", x"FFA7", x"FF9A", x"FF9A", x"FF92", x"FF9A", x"FF9C", x"FF9E", x"FFA7", x"FFA0", x"FFA6", x"FFA5", x"FFA5", x"FFAC", x"FFB1", x"FFB7", x"FFC2", x"FFC5", x"FFD1", x"FFD7", x"FFDA", x"FFDE", x"FFD4", x"FFCD", x"FFC2", x"FFBE", x"FFBF", x"FFBE", x"FFC6", x"FFC9", x"FFCA", x"FFCA", x"FFC9", x"FFC9", x"FFC5", x"FFC1", x"FFBE", x"FFBB", x"FFB9", x"FFBA", x"FFC0", x"FFC1", x"FFCC", x"FFD3", x"FFD7", x"FFDC", x"FFD8", x"FFD2", x"FFC8", x"FFC6", x"FFC7", x"FFCD", x"FFD5", x"FFE0", x"FFE4", x"FFEB", x"FFEE", x"FFF0", x"FFF4", x"FFFA", x"0001", x"000C", x"0010", x"001E", x"0020", x"0028", x"0026", x"0027", x"001E", x"0019", x"000D", x"0007", x"0002", x"0002", x"0002", x"0007", x"0007", x"0006", x"0007", x"0001", x"FFFC", x"FFF9", x"FFF0", x"FFF2", x"FFEE", x"FFF8", x"FFF9", x"FFFF", x"0001", x"0001", x"FFFF", x"0001", x"FFF6", x"FFF1", x"FFE9", x"FFE1", x"FFEA", x"FFEC", x"0000", x"0005", x"0016", x"0016", x"0020", x"001E", x"0021", x"0022", x"0024", x"0028", x"0031", x"0038", x"0043", x"004A", x"004F", x"0050", x"004C", x"0049", x"0044", x"0045", x"0045", x"0049", x"004C", x"004E", x"0049", x"004D", x"0040", x"0047", x"0035", x"0034", x"002A", x"001F", x"0022", x"0020", x"0022", x"002D", x"0030", x"003B", x"003C", x"0042", x"003F", x"003D", x"003C", x"003D", x"0044", x"004F", x"0058", x"005E", x"0067", x"006A", x"0071", x"0072", x"007D", x"0080", x"008E", x"0091", x"00A1", x"009F", x"00AE", x"00AF", x"00B4", x"00B5", x"00AD", x"00AA", x"009F", x"00A1", x"009D", x"00A3", x"00A0", x"00A4", x"00A1", x"00A0", x"009A", x"0094", x"0087", x"0087", x"0079", x"007F", x"007C", x"0084", x"0084", x"008F", x"0090", x"0095", x"0091", x"008E", x"0082", x"006F", x"0066", x"0057", x"0055", x"0056", x"0056", x"005E", x"005E", x"005C", x"005D", x"0058", x"005B", x"005E", x"0060", x"0069", x"0069", x"0076", x"0077", x"007E", x"007C", x"007B", x"0070", x"0068", x"0063", x"005D", x"005C", x"005A", x"005E", x"005D", x"005D", x"005D", x"005C", x"0057", x"0059", x"0052", x"0054", x"0056", x"005C", x"0067", x"0070", x"007F", x"0085", x"008F", x"0090", x"0091", x"0092", x"008A", x"0090", x"008A", x"0095", x"009D", x"00A5", x"00B4", x"00B4", x"00BD", x"00BA", x"00BA", x"00BA", x"00BC", x"00BE", x"00C4", x"00C7", x"00CD", x"00D3", x"00CE", x"00CF", x"00C5", x"00BF", x"00B5", x"00B5", x"00AF", x"00B3", x"00B3", x"00B6", x"00B9", x"00B8", x"00B9", x"00B5", x"00B3", x"00AD", x"00A9", x"00A3", x"009C", x"00A0", x"009F", x"00A7", x"00AA", x"00AE", x"00AB", x"00AD", x"00A2", x"009E", x"0091", x"008D", x"0082", x"0089", x"0089", x"008F", x"0093", x"009C", x"009F", x"00A6", x"00A7", x"00B1", x"00B2", x"00BB", x"00C5", x"00D0", x"00DD", x"00E8", x"00F0", x"00F2", x"00F6", x"00F0", x"00F2", x"00EB", x"00ED", x"00E9", x"00E8", x"00E9", x"00DE", x"00E3", x"00D4", x"00D0", x"00C1", x"00B7", x"00A8", x"00A4", x"009E", x"00A4", x"00A1", x"00A9", x"00A9", x"00B3", x"00B4", x"00B9", x"00B3", x"00AB", x"00A7", x"00A1", x"00A5", x"00A4", x"00B1", x"00AC", x"00BA", x"00B2", x"00B4", x"00A7", x"00A8", x"00A1", x"00A5", x"00A6", x"00AA", x"00B0", x"00B3", x"00B6", x"00B9", x"00B6", x"00BA", x"00AD", x"00B4", x"00AC", x"00AF", x"00AC", x"00B0", x"00AB", x"00AB", x"00A9", x"00AA", x"00A1", x"00A4", x"009A", x"009E", x"009C", x"00A9", x"00AE", x"00B6", x"00BD", x"00C1", x"00C3", x"00C3", x"00BC", x"00B6", x"00A8", x"00A1", x"0099", x"0092", x"0097", x"0095", x"009E", x"00A1", x"00A6", x"00A5", x"00A5", x"00A9", x"00A6", x"00B2", x"00B0", x"00BD", x"00BB", x"00CB", x"00CA", x"00C9", x"00C9", x"00B8", x"00B6", x"00AC", x"00AB", x"00A7", x"00A8", x"00A7", x"00A7", x"00A6", x"00A9", x"00A4", x"009F", x"0095", x"008F", x"0082", x"007B", x"007B", x"0077", x"007E", x"0081", x"0088", x"0088", x"008E", x"008A", x"0083", x"0083", x"0075", x"007A", x"0073", x"007E", x"007F", x"0089", x"008A", x"008C", x"0086", x"0088", x"0084", x"0086", x"008C", x"008A", x"0096", x"0094", x"009C", x"009B", x"0098", x"0097", x"008F", x"008F", x"0084", x"0088", x"007E", x"008A", x"0083", x"008B", x"0084", x"0084", x"007C", x"0072", x"006D", x"005F", x"0058", x"0055", x"0053", x"0051", x"0055", x"0052", x"0050", x"0052", x"004B", x"004A", x"003C", x"0035", x"002E", x"002B", x"0033", x"0039", x"0042", x"0049", x"004D", x"0055", x"0051", x"0054", x"0051", x"0052", x"0053", x"0058", x"0056", x"005D", x"005C", x"005B", x"0058", x"0050", x"004F", x"0045", x"004B", x"0042", x"004B", x"0047", x"004C", x"0045", x"0045", x"003E", x"0039", x"002D", x"0026", x"0014", x"000E", x"000B", x"000B", x"0014", x"0017", x"0022", x"0024", x"002D", x"002E", x"002F", x"002A", x"002B", x"0025", x"002A", x"002C", x"0031", x"0035", x"003C", x"0037", x"003D", x"0033", x"003E", x"0037", x"0040", x"0044", x"0046", x"004E", x"0052", x"0057", x"0059", x"0059", x"004E", x"004E", x"0040", x"0049", x"0040", x"004A", x"0045", x"0047", x"0044", x"0048", x"0042", x"0043", x"003A", x"0034", x"002B", x"0026", x"0029", x"0029", x"002E", x"0031", x"0035", x"0030", x"002F", x"0025", x"0016", x"0009", x"FFF9", x"FFEA", x"FFE5", x"FFE0", x"FFDF", x"FFE4", x"FFE4", x"FFE5", x"FFDF", x"FFDC", x"FFD8", x"FFDA", x"FFD6", x"FFE2", x"FFD6", x"FFE4", x"FFDF", x"FFE7", x"FFE1", x"FFE6", x"FFDA", x"FFD8", x"FFD0", x"FFCE", x"FFCC", x"FFCC", x"FFCE", x"FFCD", x"FFCE", x"FFCD", x"FFC8", x"FFC7", x"FFC3", x"FFC0", x"FFBA", x"FFBE", x"FFBB", x"FFC7", x"FFC8", x"FFD9", x"FFD4", x"FFE1", x"FFDB", x"FFDA", x"FFD8", x"FFD0", x"FFD2", x"FFCF", x"FFD5", x"FFD8", x"FFE1", x"FFE3", x"FFEC", x"FFEB", x"FFED", x"FFED", x"FFEA", x"FFEC", x"FFEB", x"FFEA", x"FFEB", x"FFE6", x"FFEB", x"FFE5", x"FFE7", x"FFE5", x"FFDB", x"FFDC", x"FFD0", x"FFD3", x"FFD0", x"FFDA", x"FFD5", x"FFD7", x"FFDA", x"FFD8", x"FFE5", x"FFED", x"FFF8", x"FFF9", x"FFF4", x"FFF6", x"FFEE", x"FFF6", x"FFF5", x"FFF6", x"FFF6", x"FFF6", x"FFF5", x"FFF8", x"FFF1", x"FFF5", x"FFF4", x"FFF2", x"FFF9", x"FFF5", x"FFF7", x"FFFB", x"FFF6", x"FFFB", x"FFF8", x"FFF9", x"FFF8", x"FFF5", x"FFF6", x"FFF7", x"FFF5", x"FFF7", x"FFF4", x"FFF6", x"FFF4", x"FFF5", x"FFF4", x"FFF4", x"FFF5", x"FFF6", x"FFF1", x"FFF8", x"FFF0", x"FFF9", x"FFF5", x"FFF6", x"FFF5", x"FFF5", x"FFF3", x"FFF3", x"FFEF", x"FFF1", x"FFEC", x"FFF0", x"FFF0", x"FFF5", x"FFF5", x"FFF9", x"FFF5", x"FFFC", x"FFF3", x"FFF8", x"FFF7", x"FFF8", x"FFFB", x"FFF8", x"FFF9", x"FFFA", x"FFF9", x"FFF7", x"FFF9", x"FFF3", x"FFF9", x"FFF6", x"FFFB", x"FFFB", x"FFFC", x"FFF9", x"FFFA", x"FFF8", x"FFFC", x"FFFB", x"FFFD", x"FFFC", x"0001", x"FFFF", x"0001", x"FFFE", x"0000", x"FFFC", x"FFFE", x"FFFA", x"FFFB", x"FFFB", x"FFFC", x"FFFA", x"FFFC", x"FFF8", x"FFFA", x"FFF5", x"FFFC", x"FFF4", x"FFFD", x"FFF6", x"FFFA", x"FFF6", x"FFF8", x"FFF6", x"FFF9", x"FFF7", x"FFF7", x"FFFB", x"FFF2", x"FFFC", x"FFF3", x"FFFB", x"FFF6", x"FFFC", x"FFF7", x"FFFF", x"FFF9", x"FFFC", x"FFFB", x"FFF7", x"FFFA", x"FFF8", x"FFFA", x"FFF6", x"FFFA", x"FFF9", x"FFF9", x"FFFB", x"FFF4", x"FFFB", x"FFF3", x"FFFA", x"FFF6", x"FFF6", x"FFF9", x"FFF5", x"FFFA", x"FFF8", x"FFF5", x"FFF9", x"FFF9", x"FFFC", x"FFFE", x"FFFC", x"0001", x"FFFC", x"0003", x"FFFE", x"0002", x"FFFF", x"FFFF", x"FFFF", x"FFFF", x"FFFE", x"FFFF", x"FFFD", x"FFFF", x"FFFD", x"FFFE", x"FFFD", x"FFFE", x"0002", x"FFFD", x"0006", x"FFFE", x"0005", x"0000", x"0002", x"0003", x"FFFF", x"0006", x"0001", x"0003", x"0007", x"FFFF", x"0005", x"0000", x"0004", x"FFFF", x"0006", x"FFFF", x"0008", x"0000", x"0009", x"0000", x"0008", x"FFFF", x"0007", x"0002", x"0004", x"0004", x"0004", x"0004", x"0006", x"0001", x"0007", x"FFFF", x"0007", x"FFFE", x"0008", x"FFFE", x"0006", x"FFFD", x"0003", x"FFFC", x"0003", x"FFFD", x"0003", x"0001", x"0001", x"0000", x"FFFC", x"0001", x"FFFB", x"0000", x"0001", x"FFFD", x"0004", x"FFFE", x"0003", x"FFFF", x"0003", x"FFFF", x"0003", x"FFFE", x"0001", x"0001", x"0001", x"0001", x"0001", x"0001", x"FFFF", x"0004", x"0001", x"0005", x"0002", x"0005", x"FFFF", x"0003", x"FFFF", x"0002", x"0002", x"0005", x"0004", x"0005", x"0006", x"0001", x"0008", x"0005", x"0007", x"0009", x"0008", x"000A", x"0008", x"000B", x"0009", x"000C", x"000B", x"0009", x"000B", x"0007", x"0009", x"0008", x"0007", x"000B", x"0007", x"000B", x"0007", x"0008", x"0008", x"0006", x"0007", x"0006", x"0003", x"0007", x"0003", x"0007", x"0005", x"0008", x"0006", x"0006", x"0006", x"0004", x"0002", x"0002", x"FFFF", x"0002", x"FFFE", x"0000", x"0000", x"FFFF", x"0002", x"FFFF", x"0002", x"0001", x"0000", x"0003", x"FFFF", x"0003", x"FFFF", x"0004", x"FFFF", x"0002", x"0000", x"0001", x"0001", x"FFFF", x"0000", x"FFFE", x"FFFD", x"0000", x"FFFD", x"FFFE", x"FFFD", x"FFFD", x"0000", x"FFFC", x"0000", x"FFFD", x"FFFF", x"FFFE", x"0002", x"FFFD", x"0003", x"FFFE", x"0001", x"0000", x"FFFF", x"0002", x"FFFD", x"0003", x"FFFE", x"0000", x"0002", x"FFFD", x"0005", x"FFFB", x"0003", x"FFFC", x"0002", x"FFFE", x"0000", x"FFFE", x"FFFF", x"FFFD", x"0000", x"FFFE", x"FFFF", x"0001", x"FFFD", x"0005", x"FFFE", x"0002", x"0003", x"0001", x"0006", x"0002", x"0007", x"0000", x"0006", x"0000", x"0003", x"0003", x"0001", x"0001", x"0005", x"0003", x"0004", x"0005", x"FFFF", x"0007", x"0000", x"0005", x"0002", x"0004", x"0000", x"0002", x"0000", x"FFFF", x"0003", x"FFFE", x"0004", x"0000", x"0002", x"0003", x"0000", x"0004", x"0002", x"FFFF", x"0003", x"0004", x"0001", x"0009", x"0000", x"0006", x"0003", x"0004", x"0005", x"0003", x"0003", x"0002", x"0005", x"0000", x"0003", x"0002", x"0004", x"0002", x"0005", x"0000", x"0006", x"0001", x"0006", x"0001", x"0003", x"0002", x"0001", x"0004", x"0000", x"0006", x"0001", x"0004", x"0001", x"0001", x"0005", x"FFFF", x"0005", x"FFFF", x"0001", x"0001", x"FFFE", x"0000", x"FFFE", x"FFFF", x"0000", x"FFFE", x"FFFF", x"0001", x"0000", x"0000", x"0000", x"0001", x"0004", x"0006", x"0005", x"0004", x"0006", x"0006", x"0006", x"0006", x"0004", x"0004", x"0004", x"0001", x"0001", x"0001", x"0001", x"FFFE", x"0001", x"FFFF", x"0003", x"FFFF", x"0001", x"0000", x"0003", x"0001", x"0003", x"0002", x"0002", x"0002", x"0002", x"0001", x"0001", x"0002", x"0001", x"FFFE", x"0005", x"FFFF", x"0003", x"0003", x"0001", x"0004", x"FFFF", x"0003", x"0001", x"0003", x"0002", x"0001", x"0001", x"0004", x"0002", x"0005", x"0000", x"0004", x"FFFF", x"0001", x"0002", x"FFFF", x"0004", x"0003", x"0002", x"0006", x"0001", x"0008", x"FFFF", x"0007", x"0001", x"0004", x"0003", x"0003", x"0000", x"0006", x"FFFF", x"0006", x"0000", x"0001", x"0002", x"FFFF", x"FFFF", x"0002", x"FFFE", x"0004", x"0001", x"0000", x"0002", x"0002", x"FFFF", x"0002", x"FFFE", x"0004", x"FFFE", x"0005", x"FFFE", x"0005", x"FFFF", x"0003", x"FFFF", x"0003", x"0001", x"0001", x"0002", x"0000", x"0004", x"0000", x"0004", x"FFFF", x"0005", x"FFFC", x"0005", x"FFFE", x"0004", x"FFFE", x"0003", x"FFFE", x"0006", x"FFFF", x"0002", x"0000", x"0001", x"0002", x"0000", x"0002", x"FFFF", x"0001", x"0002", x"0000", x"0002", x"0003", x"0000", x"0003", x"FFFF", x"0003", x"FFFF", x"0004", x"FFFF", x"0001", x"0000", x"FFFE", x"0001", x"FFFC", x"0002", x"FFFC", x"0003", x"FFFC", x"0005", x"FFFB", x"0006", x"FFFC", x"0002", x"0002", x"0001", x"0003", x"0000", x"0003", x"0001", x"0003", x"0001", x"0003", x"FFFF", x"0001", x"0000", x"0000", x"0001", x"0001", x"0001", x"FFFE", x"0002", x"FFFF", x"0000", x"0003", x"FFFE", x"0002", x"FFFF", x"0000", x"0002", x"0000", x"0004", x"FFFF", x"0004", x"FFFE", x"0003", x"0000", x"0001", x"0000", x"0000", x"0001", x"0002", x"FFFF", x"0004", x"FFFF", x"0003", x"0000", x"0001", x"0002", x"FFFF", x"0003", x"0000", x"0000", x"0000", x"0001", x"FFFE", x"0003", x"FFFF", x"0003", x"FFFF", x"0003", x"FFFF", x"0003", x"0000", x"0002", x"0001", x"0003", x"0000", x"0005", x"FFFF", x"0004", x"0002", x"0000", x"0002", x"0001", x"0001", x"0004", x"0002", x"0001", x"0002", x"FFFF", x"0004", x"FFFE", x"0006", x"FFFE", x"0004", x"FFFE", x"0005", x"FFFB", x"0008", x"FFFA", x"0004", x"FFFE", x"0000", x"0002", x"FFFD", x"0004", x"FFFB", x"0007", x"FFFF", x"0007", x"0003", x"0004", x"0004", x"0004", x"0001", x"0005", x"0001", x"0005", x"0001", x"0005", x"0000", x"0002", x"0003", x"0000", x"0004", x"0002", x"0000", x"0002", x"0000", x"0004", x"0001", x"0004", x"0004", x"0003", x"0005", x"0000", x"0005", x"0000", x"0002", x"0004", x"FFFF", x"0005", x"FFFF", x"0003", x"0001", x"0002", x"0004", x"FFFE", x"0005", x"FFFE", x"0005", x"0001", x"0002", x"0000", x"0002", x"0001", x"0000", x"0003", x"FFFE", x"0004", x"FFFC", x"0003", x"FFFE", x"0001", x"0003", x"FFFF", x"0002", x"0000", x"0002", x"FFFF", x"0002", x"0000", x"0002", x"0000", x"0002", x"0000", x"0003", x"0001", x"0002", x"0003", x"FFFE", x"0003", x"FFFD", x"0004", x"FFFE", x"0003", x"FFFD", x"0003", x"FFFE", x"0001", x"0001", x"FFFF", x"0000", x"FFFF", x"0002", x"FFFF", x"0004", x"0002", x"0003", x"0004", x"0001", x"0003", x"0001", x"0003", x"0002", x"0002", x"0003", x"0003", x"0003", x"0003", x"0003", x"0001", x"0002", x"0003", x"0000", x"0004", x"0000", x"0004", x"0002", x"0004", x"0001", x"0003", x"0004", x"0001", x"0004", x"FFFE", x"0004", x"FFFC", x"0002", x"FFFF", x"0000", x"0002", x"FFFF", x"0003", x"FFFF", x"0003", x"0000", x"0001", x"0002", x"0001", x"0001", x"FFFF", x"0003", x"FFFF", x"0003", x"FFFF", x"0002", x"FFFE", x"0002", x"0001", x"0001", x"0003", x"FFFF", x"0003", x"0001", x"0002", x"0000", x"0002", x"0002", x"FFFF", x"0001", x"0002", x"FFFF", x"0006", x"FFFE", x"0006", x"FFFC", x"0005", x"FFFF", x"0000", x"0001", x"FFFE", x"0001", x"FFFF", x"FFFE", x"0003", x"FFFE", x"0004", x"FFFF", x"0003", x"FFFF", x"0001", x"FFFE", x"FFFF", x"0001", x"FFFF", x"0005", x"FFFE", x"0003", x"0000", x"0003", x"0002", x"0002", x"0001", x"0003", x"0000", x"0003", x"0002", x"0000", x"0003", x"FFFD", x"0006", x"FFFD", x"0004", x"FFFF", x"0001", x"0004", x"FFFF", x"0001", x"0000", x"0000", x"0002", x"0000", x"0005", x"0001", x"0003", x"FFFF", x"0002", x"0000", x"0003", x"0001", x"0001", x"0004", x"FFFD", x"0004", x"0000", x"FFFF", x"0001", x"0001", x"0000", x"0001", x"0000", x"FFFE", x"0001", x"0000", x"0004", x"0000", x"0002", x"FFFF", x"0000", x"0000", x"0002", x"0001", x"0004", x"0000", x"0002", x"0001", x"0000", x"0002", x"0000", x"0003", x"0001", x"0003", x"0000", x"0004", x"FFFF", x"0004", x"FFFE", x"0003", x"0000", x"0001", x"0001", x"FFFF", x"0000", x"0002", x"FFFF", x"0001", x"FFFF", x"0001", x"FFFF", x"0001", x"FFFD", x"0001", x"FFFD", x"0001", x"0000", x"FFFF", x"0002", x"FFFE", x"0003", x"FFFF", x"FFFF", x"0002", x"FFFE", x"0001", x"0001", x"FFFE", x"0002", x"FFFF", x"FFFF", x"0001", x"FFFF", x"FFFD", x"0002", x"FFF8", x"0001", x"FFFB", x"FFFD", x"0001", x"FFFE", x"0001", x"0000", x"0000", x"FFFD", x"0002", x"FFFC", x"0002", x"FFFD", x"FFFF", x"0000", x"0000", x"0001", x"FFFF", x"0001", x"FFFF", x"0002", x"FFFE", x"FFFF", x"FFFE", x"FFFE", x"FFFE", x"0002", x"FFFD", x"0003", x"FFFD", x"0003", x"FFFE", x"0002", x"0001", x"0000", x"0001", x"0001", x"0000", x"0002", x"0001", x"FFFE", x"0000", x"FFFD", x"FFFF", x"0000", x"FFFD", x"0002", x"FFFB", x"0004", x"FFFE", x"0003", x"0000", x"0001", x"0001", x"0003", x"FFFD", x"0004", x"FFFC", x"0003", x"FFFE", x"FFFD", x"0000", x"FFFF", x"FFFF", x"0002", x"0000", x"FFFF", x"0002", x"FFFE", x"FFFF", x"0001", x"FFFC", x"0003", x"FFFA", x"0004", x"FFF9", x"0004", x"FFFA", x"0006", x"FFFA", x"0006", x"FFFB", x"0002", x"0001", x"FFFD", x"0004", x"FFFD", x"0001", x"FFFF", x"0000", x"FFFE", x"0000", x"FFFE", x"0000", x"0002", x"FFFE", x"0002", x"FFFE", x"0000", x"FFFF", x"FFFF", x"0001", x"FFFD", x"0001", x"FFFD", x"FFFF", x"FFFF", x"FFFE", x"0001", x"FFF9", x"0004", x"FFFB", x"0001", x"FFFF", x"FFFD", x"FFFD", x"0000", x"FFFB", x"0001", x"FFFD", x"0000", x"FFFF", x"FFFE", x"0001", x"0000", x"0000", x"0002", x"FFFF", x"0002", x"0000", x"0002", x"FFFF", x"0000", x"0001", x"FFFF", x"FFFF", x"FFFF", x"FFFC", x"0000", x"FFFB", x"0003", x"FFFB", x"0004", x"FFFE", x"0001", x"0000", x"0002", x"0000", x"FFFF", x"0001", x"FFFB", x"0000", x"FFFC", x"0000", x"FFFC", x"0002", x"FFFC", x"0002", x"FFFD", x"0003", x"FFFD", x"0001", x"FFFF", x"FFFF", x"FFFF", x"FFFE", x"0001", x"FFFC", x"0005", x"FFFA", x"0003", x"FFFC", x"FFFF", x"0001", x"FFFB", x"0003", x"FFFC", x"0000", x"FFFE", x"FFFF", x"FFFF", x"0000", x"0001", x"FFFD", x"FFFF", x"FFFE", x"FFFE", x"FFFF", x"FFFE", x"0000", x"FFFE", x"0000", x"FFFD", x"FFFD", x"FFFF", x"FFF9", x"FFFF", x"FFFB", x"FFFF", x"FFFE", x"FFFF", x"FFFF", x"FFFE", x"FFFE", x"FFFF", x"FFFF", x"0001", x"FFFF", x"0000", x"FFFD", x"0001", x"FFFE", x"0003", x"FFFF", x"0002", x"FFFE", x"0002", x"FFFF", x"0000", x"0001", x"FFFF", x"0003", x"FFFD", x"0003", x"FFFD", x"0002", x"FFFF", x"0001", x"0001", x"FFFE", x"0001", x"FFFB", x"0002", x"FFFA", x"0001", x"FFFF", x"FFFE", x"0001", x"FFFD", x"0001", x"FFFF", x"0001", x"FFFE", x"FFFE", x"FFFE", x"FFFF", x"FFFD", x"0002", x"FFFE", x"FFFF", x"0000", x"FFFD", x"0001", x"FFFD", x"0001", x"FFFC", x"FFFD", x"FFFE", x"FFFC", x"0002", x"FFFB", x"0004", x"FFFC", x"0003", x"FFFE", x"0002", x"FFFD", x"0006", x"FFFC", x"0004", x"0000", x"0001", x"0001", x"0002", x"FFFE", x"0005", x"FFFD", x"0003", x"FFFC", x"0000", x"0000", x"FFFC", x"0001", x"FFFE", x"FFFF", x"0000", x"FFFE", x"0002", x"FFFE", x"0005", x"FFFA", x"0004", x"FFFB", x"0002", x"FFFE", x"FFFF", x"FFFE", x"FFFD", x"FFFE", x"FFFB", x"0000", x"FFFA", x"0001", x"FFFC", x"FFFF", x"FFFF", x"FFFE", x"0001", x"FFFE", x"0001", x"0000", x"FFFC", x"0003", x"FFFB", x"0002", x"FFFE", x"FFFF", x"FFFE", x"0002", x"FFFD", x"0005", x"FFFA", x"0005", x"FFF9", x"0003", x"FFFB", x"0003", x"FFFC", x"0002", x"0000");
--  constant SoundR : TROM := (x"0000", x"30FB", x"5A82", x"7641", x"7FFF", x"7641", x"5A82", x"30FB", x"0000", x"CF05", x"A57E", x"89BF", x"8001", x"89BF", x"A57E", x"CF05");
  signal Counter : natural := 0;
begin
  process(iClk)
  begin
    if(rising_edge(iClk)) then
      if(iRst = '1') then
        Counter <= 0;
      elsif(iEn = '1') then
        if(Counter < ArraySize) then
          Counter <= Counter + 1;
        else
          Counter <= 0;
        end if;
      end if;
    end if;
  end process;
  oDataL <= SoundL(Counter);
  oDataR <= SoundL(Counter);
end RTL;